initial begin
RAM[16'h0000] = 8'h00;
RAM[16'h0001] = 8'h00;
RAM[16'h0002] = 8'h00;
RAM[16'h0003] = 8'h00;
RAM[16'h0004] = 8'h00;
RAM[16'h0005] = 8'h00;
RAM[16'h0006] = 8'h00;
RAM[16'h0007] = 8'h00;
RAM[16'h0008] = 8'h00;
RAM[16'h0009] = 8'h00;
RAM[16'h000A] = 8'h00;
RAM[16'h000B] = 8'h00;
RAM[16'h000C] = 8'h00;
RAM[16'h000D] = 8'h00;
RAM[16'h000E] = 8'h00;
RAM[16'h000F] = 8'h00;
RAM[16'h0010] = 8'h00;
RAM[16'h0011] = 8'h00;
RAM[16'h0012] = 8'h00;
RAM[16'h0013] = 8'h00;
RAM[16'h0014] = 8'h00;
RAM[16'h0015] = 8'h00;
RAM[16'h0016] = 8'h00;
RAM[16'h0017] = 8'h00;
RAM[16'h0018] = 8'h00;
RAM[16'h0019] = 8'h00;
RAM[16'h001A] = 8'h00;
RAM[16'h001B] = 8'h00;
RAM[16'h001C] = 8'h00;
RAM[16'h001D] = 8'h00;
RAM[16'h001E] = 8'h00;
RAM[16'h001F] = 8'h00;
RAM[16'h0020] = 8'h00;
RAM[16'h0021] = 8'h00;
RAM[16'h0022] = 8'h00;
RAM[16'h0023] = 8'h00;
RAM[16'h0024] = 8'h00;
RAM[16'h0025] = 8'h00;
RAM[16'h0026] = 8'h00;
RAM[16'h0027] = 8'h00;
RAM[16'h0028] = 8'h00;
RAM[16'h0029] = 8'h00;
RAM[16'h002A] = 8'h00;
RAM[16'h002B] = 8'h00;
RAM[16'h002C] = 8'h00;
RAM[16'h002D] = 8'h00;
RAM[16'h002E] = 8'h00;
RAM[16'h002F] = 8'h00;
RAM[16'h0030] = 8'h00;
RAM[16'h0031] = 8'h00;
RAM[16'h0032] = 8'h00;
RAM[16'h0033] = 8'h00;
RAM[16'h0034] = 8'h00;
RAM[16'h0035] = 8'h00;
RAM[16'h0036] = 8'h00;
RAM[16'h0037] = 8'h00;
RAM[16'h0038] = 8'h00;
RAM[16'h0039] = 8'h00;
RAM[16'h003A] = 8'h00;
RAM[16'h003B] = 8'h00;
RAM[16'h003C] = 8'h00;
RAM[16'h003D] = 8'h00;
RAM[16'h003E] = 8'h00;
RAM[16'h003F] = 8'h00;
RAM[16'h0040] = 8'h00;
RAM[16'h0041] = 8'h00;
RAM[16'h0042] = 8'h00;
RAM[16'h0043] = 8'h00;
RAM[16'h0044] = 8'h00;
RAM[16'h0045] = 8'h00;
RAM[16'h0046] = 8'h00;
RAM[16'h0047] = 8'h00;
RAM[16'h0048] = 8'h00;
RAM[16'h0049] = 8'h00;
RAM[16'h004A] = 8'h00;
RAM[16'h004B] = 8'h00;
RAM[16'h004C] = 8'h00;
RAM[16'h004D] = 8'h00;
RAM[16'h004E] = 8'h00;
RAM[16'h004F] = 8'h00;
RAM[16'h0050] = 8'h00;
RAM[16'h0051] = 8'h00;
RAM[16'h0052] = 8'h00;
RAM[16'h0053] = 8'h00;
RAM[16'h0054] = 8'h00;
RAM[16'h0055] = 8'h00;
RAM[16'h0056] = 8'h00;
RAM[16'h0057] = 8'h00;
RAM[16'h0058] = 8'h00;
RAM[16'h0059] = 8'h00;
RAM[16'h005A] = 8'h00;
RAM[16'h005B] = 8'h00;
RAM[16'h005C] = 8'h00;
RAM[16'h005D] = 8'h00;
RAM[16'h005E] = 8'h00;
RAM[16'h005F] = 8'h00;
RAM[16'h0060] = 8'h00;
RAM[16'h0061] = 8'h00;
RAM[16'h0062] = 8'h00;
RAM[16'h0063] = 8'h00;
RAM[16'h0064] = 8'h00;
RAM[16'h0065] = 8'h00;
RAM[16'h0066] = 8'h00;
RAM[16'h0067] = 8'h00;
RAM[16'h0068] = 8'h00;
RAM[16'h0069] = 8'h00;
RAM[16'h006A] = 8'h00;
RAM[16'h006B] = 8'h00;
RAM[16'h006C] = 8'h00;
RAM[16'h006D] = 8'h00;
RAM[16'h006E] = 8'h00;
RAM[16'h006F] = 8'h00;
RAM[16'h0070] = 8'h00;
RAM[16'h0071] = 8'h00;
RAM[16'h0072] = 8'h00;
RAM[16'h0073] = 8'h00;
RAM[16'h0074] = 8'h00;
RAM[16'h0075] = 8'h00;
RAM[16'h0076] = 8'h00;
RAM[16'h0077] = 8'h00;
RAM[16'h0078] = 8'h00;
RAM[16'h0079] = 8'h00;
RAM[16'h007A] = 8'h00;
RAM[16'h007B] = 8'h00;
RAM[16'h007C] = 8'h00;
RAM[16'h007D] = 8'h00;
RAM[16'h007E] = 8'h00;
RAM[16'h007F] = 8'h00;
RAM[16'h0080] = 8'h00;
RAM[16'h0081] = 8'h00;
RAM[16'h0082] = 8'h00;
RAM[16'h0083] = 8'h00;
RAM[16'h0084] = 8'h00;
RAM[16'h0085] = 8'h00;
RAM[16'h0086] = 8'h00;
RAM[16'h0087] = 8'h00;
RAM[16'h0088] = 8'h00;
RAM[16'h0089] = 8'h00;
RAM[16'h008A] = 8'h00;
RAM[16'h008B] = 8'h00;
RAM[16'h008C] = 8'h00;
RAM[16'h008D] = 8'h00;
RAM[16'h008E] = 8'h00;
RAM[16'h008F] = 8'h00;
RAM[16'h0090] = 8'h00;
RAM[16'h0091] = 8'h00;
RAM[16'h0092] = 8'h00;
RAM[16'h0093] = 8'h00;
RAM[16'h0094] = 8'h00;
RAM[16'h0095] = 8'h00;
RAM[16'h0096] = 8'h00;
RAM[16'h0097] = 8'h00;
RAM[16'h0098] = 8'h00;
RAM[16'h0099] = 8'h00;
RAM[16'h009A] = 8'h00;
RAM[16'h009B] = 8'h00;
RAM[16'h009C] = 8'h00;
RAM[16'h009D] = 8'h00;
RAM[16'h009E] = 8'h00;
RAM[16'h009F] = 8'h00;
RAM[16'h00A0] = 8'h00;
RAM[16'h00A1] = 8'h00;
RAM[16'h00A2] = 8'h00;
RAM[16'h00A3] = 8'h00;
RAM[16'h00A4] = 8'h00;
RAM[16'h00A5] = 8'h00;
RAM[16'h00A6] = 8'h00;
RAM[16'h00A7] = 8'h00;
RAM[16'h00A8] = 8'h00;
RAM[16'h00A9] = 8'h00;
RAM[16'h00AA] = 8'h00;
RAM[16'h00AB] = 8'h00;
RAM[16'h00AC] = 8'h00;
RAM[16'h00AD] = 8'h00;
RAM[16'h00AE] = 8'h00;
RAM[16'h00AF] = 8'h00;
RAM[16'h00B0] = 8'h00;
RAM[16'h00B1] = 8'h00;
RAM[16'h00B2] = 8'h00;
RAM[16'h00B3] = 8'h00;
RAM[16'h00B4] = 8'h00;
RAM[16'h00B5] = 8'h00;
RAM[16'h00B6] = 8'h00;
RAM[16'h00B7] = 8'h00;
RAM[16'h00B8] = 8'h00;
RAM[16'h00B9] = 8'h00;
RAM[16'h00BA] = 8'h00;
RAM[16'h00BB] = 8'h00;
RAM[16'h00BC] = 8'h00;
RAM[16'h00BD] = 8'h00;
RAM[16'h00BE] = 8'h00;
RAM[16'h00BF] = 8'h00;
RAM[16'h00C0] = 8'h00;
RAM[16'h00C1] = 8'h00;
RAM[16'h00C2] = 8'h00;
RAM[16'h00C3] = 8'h00;
RAM[16'h00C4] = 8'h00;
RAM[16'h00C5] = 8'h00;
RAM[16'h00C6] = 8'h00;
RAM[16'h00C7] = 8'h00;
RAM[16'h00C8] = 8'h00;
RAM[16'h00C9] = 8'h00;
RAM[16'h00CA] = 8'h00;
RAM[16'h00CB] = 8'h00;
RAM[16'h00CC] = 8'h00;
RAM[16'h00CD] = 8'h00;
RAM[16'h00CE] = 8'h00;
RAM[16'h00CF] = 8'h00;
RAM[16'h00D0] = 8'h00;
RAM[16'h00D1] = 8'h00;
RAM[16'h00D2] = 8'h00;
RAM[16'h00D3] = 8'h00;
RAM[16'h00D4] = 8'h00;
RAM[16'h00D5] = 8'h00;
RAM[16'h00D6] = 8'h00;
RAM[16'h00D7] = 8'h00;
RAM[16'h00D8] = 8'h00;
RAM[16'h00D9] = 8'h00;
RAM[16'h00DA] = 8'h00;
RAM[16'h00DB] = 8'h00;
RAM[16'h00DC] = 8'h00;
RAM[16'h00DD] = 8'h00;
RAM[16'h00DE] = 8'h00;
RAM[16'h00DF] = 8'h00;
RAM[16'h00E0] = 8'h00;
RAM[16'h00E1] = 8'h00;
RAM[16'h00E2] = 8'h00;
RAM[16'h00E3] = 8'h00;
RAM[16'h00E4] = 8'h00;
RAM[16'h00E5] = 8'h00;
RAM[16'h00E6] = 8'h00;
RAM[16'h00E7] = 8'h00;
RAM[16'h00E8] = 8'h00;
RAM[16'h00E9] = 8'h00;
RAM[16'h00EA] = 8'h00;
RAM[16'h00EB] = 8'h00;
RAM[16'h00EC] = 8'h00;
RAM[16'h00ED] = 8'h00;
RAM[16'h00EE] = 8'h00;
RAM[16'h00EF] = 8'h00;
RAM[16'h00F0] = 8'h00;
RAM[16'h00F1] = 8'h00;
RAM[16'h00F2] = 8'h00;
RAM[16'h00F3] = 8'h00;
RAM[16'h00F4] = 8'h00;
RAM[16'h00F5] = 8'h00;
RAM[16'h00F6] = 8'h00;
RAM[16'h00F7] = 8'h00;
RAM[16'h00F8] = 8'h00;
RAM[16'h00F9] = 8'h00;
RAM[16'h00FA] = 8'h00;
RAM[16'h00FB] = 8'h00;
RAM[16'h00FC] = 8'h00;
RAM[16'h00FD] = 8'h00;
RAM[16'h00FE] = 8'h00;
RAM[16'h00FF] = 8'h00;
RAM[16'h0100] = 8'h00;
RAM[16'h0101] = 8'h00;
RAM[16'h0102] = 8'h00;
RAM[16'h0103] = 8'h00;
RAM[16'h0104] = 8'h00;
RAM[16'h0105] = 8'h00;
RAM[16'h0106] = 8'h00;
RAM[16'h0107] = 8'h00;
RAM[16'h0108] = 8'h00;
RAM[16'h0109] = 8'h00;
RAM[16'h010A] = 8'h00;
RAM[16'h010B] = 8'h00;
RAM[16'h010C] = 8'h00;
RAM[16'h010D] = 8'h00;
RAM[16'h010E] = 8'h00;
RAM[16'h010F] = 8'h00;
RAM[16'h0110] = 8'h00;
RAM[16'h0111] = 8'h00;
RAM[16'h0112] = 8'h00;
RAM[16'h0113] = 8'h00;
RAM[16'h0114] = 8'h00;
RAM[16'h0115] = 8'h00;
RAM[16'h0116] = 8'h00;
RAM[16'h0117] = 8'h00;
RAM[16'h0118] = 8'h00;
RAM[16'h0119] = 8'h00;
RAM[16'h011A] = 8'h00;
RAM[16'h011B] = 8'h00;
RAM[16'h011C] = 8'h00;
RAM[16'h011D] = 8'h00;
RAM[16'h011E] = 8'h00;
RAM[16'h011F] = 8'h00;
RAM[16'h0120] = 8'h00;
RAM[16'h0121] = 8'h00;
RAM[16'h0122] = 8'h00;
RAM[16'h0123] = 8'h00;
RAM[16'h0124] = 8'h00;
RAM[16'h0125] = 8'h00;
RAM[16'h0126] = 8'h00;
RAM[16'h0127] = 8'h00;
RAM[16'h0128] = 8'h00;
RAM[16'h0129] = 8'h00;
RAM[16'h012A] = 8'h00;
RAM[16'h012B] = 8'h00;
RAM[16'h012C] = 8'h00;
RAM[16'h012D] = 8'h00;
RAM[16'h012E] = 8'h00;
RAM[16'h012F] = 8'h00;
RAM[16'h0130] = 8'h00;
RAM[16'h0131] = 8'h00;
RAM[16'h0132] = 8'h00;
RAM[16'h0133] = 8'h00;
RAM[16'h0134] = 8'h00;
RAM[16'h0135] = 8'h00;
RAM[16'h0136] = 8'h00;
RAM[16'h0137] = 8'h00;
RAM[16'h0138] = 8'h00;
RAM[16'h0139] = 8'h00;
RAM[16'h013A] = 8'h00;
RAM[16'h013B] = 8'h00;
RAM[16'h013C] = 8'h00;
RAM[16'h013D] = 8'h00;
RAM[16'h013E] = 8'h00;
RAM[16'h013F] = 8'h00;
RAM[16'h0140] = 8'h00;
RAM[16'h0141] = 8'h00;
RAM[16'h0142] = 8'h00;
RAM[16'h0143] = 8'h00;
RAM[16'h0144] = 8'h00;
RAM[16'h0145] = 8'h00;
RAM[16'h0146] = 8'h00;
RAM[16'h0147] = 8'h00;
RAM[16'h0148] = 8'h00;
RAM[16'h0149] = 8'h00;
RAM[16'h014A] = 8'h00;
RAM[16'h014B] = 8'h00;
RAM[16'h014C] = 8'h00;
RAM[16'h014D] = 8'h00;
RAM[16'h014E] = 8'h00;
RAM[16'h014F] = 8'h00;
RAM[16'h0150] = 8'h00;
RAM[16'h0151] = 8'h00;
RAM[16'h0152] = 8'h00;
RAM[16'h0153] = 8'h00;
RAM[16'h0154] = 8'h00;
RAM[16'h0155] = 8'h00;
RAM[16'h0156] = 8'h00;
RAM[16'h0157] = 8'h00;
RAM[16'h0158] = 8'h00;
RAM[16'h0159] = 8'h00;
RAM[16'h015A] = 8'h00;
RAM[16'h015B] = 8'h00;
RAM[16'h015C] = 8'h00;
RAM[16'h015D] = 8'h00;
RAM[16'h015E] = 8'h00;
RAM[16'h015F] = 8'h00;
RAM[16'h0160] = 8'h00;
RAM[16'h0161] = 8'h00;
RAM[16'h0162] = 8'h00;
RAM[16'h0163] = 8'h00;
RAM[16'h0164] = 8'h00;
RAM[16'h0165] = 8'h00;
RAM[16'h0166] = 8'h00;
RAM[16'h0167] = 8'h00;
RAM[16'h0168] = 8'h00;
RAM[16'h0169] = 8'h00;
RAM[16'h016A] = 8'h00;
RAM[16'h016B] = 8'h00;
RAM[16'h016C] = 8'h00;
RAM[16'h016D] = 8'h00;
RAM[16'h016E] = 8'h00;
RAM[16'h016F] = 8'h00;
RAM[16'h0170] = 8'h00;
RAM[16'h0171] = 8'h00;
RAM[16'h0172] = 8'h00;
RAM[16'h0173] = 8'h00;
RAM[16'h0174] = 8'h00;
RAM[16'h0175] = 8'h00;
RAM[16'h0176] = 8'h00;
RAM[16'h0177] = 8'h00;
RAM[16'h0178] = 8'h00;
RAM[16'h0179] = 8'h00;
RAM[16'h017A] = 8'h00;
RAM[16'h017B] = 8'h00;
RAM[16'h017C] = 8'h00;
RAM[16'h017D] = 8'h00;
RAM[16'h017E] = 8'h00;
RAM[16'h017F] = 8'h00;
RAM[16'h0180] = 8'h00;
RAM[16'h0181] = 8'h00;
RAM[16'h0182] = 8'h00;
RAM[16'h0183] = 8'h00;
RAM[16'h0184] = 8'h00;
RAM[16'h0185] = 8'h00;
RAM[16'h0186] = 8'h00;
RAM[16'h0187] = 8'h00;
RAM[16'h0188] = 8'h00;
RAM[16'h0189] = 8'h00;
RAM[16'h018A] = 8'h00;
RAM[16'h018B] = 8'h00;
RAM[16'h018C] = 8'h00;
RAM[16'h018D] = 8'h00;
RAM[16'h018E] = 8'h00;
RAM[16'h018F] = 8'h00;
RAM[16'h0190] = 8'h00;
RAM[16'h0191] = 8'h00;
RAM[16'h0192] = 8'h00;
RAM[16'h0193] = 8'h00;
RAM[16'h0194] = 8'h00;
RAM[16'h0195] = 8'h00;
RAM[16'h0196] = 8'h00;
RAM[16'h0197] = 8'h00;
RAM[16'h0198] = 8'h00;
RAM[16'h0199] = 8'h00;
RAM[16'h019A] = 8'h00;
RAM[16'h019B] = 8'h00;
RAM[16'h019C] = 8'h00;
RAM[16'h019D] = 8'h00;
RAM[16'h019E] = 8'h00;
RAM[16'h019F] = 8'h00;
RAM[16'h01A0] = 8'h00;
RAM[16'h01A1] = 8'h00;
RAM[16'h01A2] = 8'h00;
RAM[16'h01A3] = 8'h00;
RAM[16'h01A4] = 8'h00;
RAM[16'h01A5] = 8'h00;
RAM[16'h01A6] = 8'h00;
RAM[16'h01A7] = 8'h00;
RAM[16'h01A8] = 8'h00;
RAM[16'h01A9] = 8'h00;
RAM[16'h01AA] = 8'h00;
RAM[16'h01AB] = 8'h00;
RAM[16'h01AC] = 8'h00;
RAM[16'h01AD] = 8'h00;
RAM[16'h01AE] = 8'h00;
RAM[16'h01AF] = 8'h00;
RAM[16'h01B0] = 8'h00;
RAM[16'h01B1] = 8'h00;
RAM[16'h01B2] = 8'h00;
RAM[16'h01B3] = 8'h00;
RAM[16'h01B4] = 8'h00;
RAM[16'h01B5] = 8'h00;
RAM[16'h01B6] = 8'h00;
RAM[16'h01B7] = 8'h00;
RAM[16'h01B8] = 8'h00;
RAM[16'h01B9] = 8'h00;
RAM[16'h01BA] = 8'h00;
RAM[16'h01BB] = 8'h00;
RAM[16'h01BC] = 8'h00;
RAM[16'h01BD] = 8'h00;
RAM[16'h01BE] = 8'h00;
RAM[16'h01BF] = 8'h00;
RAM[16'h01C0] = 8'h00;
RAM[16'h01C1] = 8'h00;
RAM[16'h01C2] = 8'h00;
RAM[16'h01C3] = 8'h00;
RAM[16'h01C4] = 8'h00;
RAM[16'h01C5] = 8'h00;
RAM[16'h01C6] = 8'h00;
RAM[16'h01C7] = 8'h00;
RAM[16'h01C8] = 8'h00;
RAM[16'h01C9] = 8'h00;
RAM[16'h01CA] = 8'h00;
RAM[16'h01CB] = 8'h00;
RAM[16'h01CC] = 8'h00;
RAM[16'h01CD] = 8'h00;
RAM[16'h01CE] = 8'h00;
RAM[16'h01CF] = 8'h00;
RAM[16'h01D0] = 8'h00;
RAM[16'h01D1] = 8'h00;
RAM[16'h01D2] = 8'h00;
RAM[16'h01D3] = 8'h00;
RAM[16'h01D4] = 8'h00;
RAM[16'h01D5] = 8'h00;
RAM[16'h01D6] = 8'h00;
RAM[16'h01D7] = 8'h00;
RAM[16'h01D8] = 8'h00;
RAM[16'h01D9] = 8'h00;
RAM[16'h01DA] = 8'h00;
RAM[16'h01DB] = 8'h00;
RAM[16'h01DC] = 8'h00;
RAM[16'h01DD] = 8'h00;
RAM[16'h01DE] = 8'h00;
RAM[16'h01DF] = 8'h00;
RAM[16'h01E0] = 8'h00;
RAM[16'h01E1] = 8'h00;
RAM[16'h01E2] = 8'h00;
RAM[16'h01E3] = 8'h00;
RAM[16'h01E4] = 8'h00;
RAM[16'h01E5] = 8'h00;
RAM[16'h01E6] = 8'h00;
RAM[16'h01E7] = 8'h00;
RAM[16'h01E8] = 8'h00;
RAM[16'h01E9] = 8'h00;
RAM[16'h01EA] = 8'h00;
RAM[16'h01EB] = 8'h00;
RAM[16'h01EC] = 8'h00;
RAM[16'h01ED] = 8'h00;
RAM[16'h01EE] = 8'h00;
RAM[16'h01EF] = 8'h00;
RAM[16'h01F0] = 8'h00;
RAM[16'h01F1] = 8'h00;
RAM[16'h01F2] = 8'h00;
RAM[16'h01F3] = 8'h00;
RAM[16'h01F4] = 8'h00;
RAM[16'h01F5] = 8'h00;
RAM[16'h01F6] = 8'h00;
RAM[16'h01F7] = 8'h00;
RAM[16'h01F8] = 8'h00;
RAM[16'h01F9] = 8'h00;
RAM[16'h01FA] = 8'h00;
RAM[16'h01FB] = 8'h00;
RAM[16'h01FC] = 8'h00;
RAM[16'h01FD] = 8'h00;
RAM[16'h01FE] = 8'h00;
RAM[16'h01FF] = 8'h00;
RAM[16'h0200] = 8'h00;
RAM[16'h0201] = 8'h00;
RAM[16'h0202] = 8'h00;
RAM[16'h0203] = 8'h00;
RAM[16'h0204] = 8'h00;
RAM[16'h0205] = 8'h00;
RAM[16'h0206] = 8'h00;
RAM[16'h0207] = 8'h00;
RAM[16'h0208] = 8'h00;
RAM[16'h0209] = 8'h00;
RAM[16'h020A] = 8'h00;
RAM[16'h020B] = 8'h00;
RAM[16'h020C] = 8'h00;
RAM[16'h020D] = 8'h00;
RAM[16'h020E] = 8'h00;
RAM[16'h020F] = 8'h00;
RAM[16'h0210] = 8'h00;
RAM[16'h0211] = 8'h00;
RAM[16'h0212] = 8'h00;
RAM[16'h0213] = 8'h00;
RAM[16'h0214] = 8'h00;
RAM[16'h0215] = 8'h00;
RAM[16'h0216] = 8'h00;
RAM[16'h0217] = 8'h00;
RAM[16'h0218] = 8'h00;
RAM[16'h0219] = 8'h00;
RAM[16'h021A] = 8'h00;
RAM[16'h021B] = 8'h00;
RAM[16'h021C] = 8'h00;
RAM[16'h021D] = 8'h00;
RAM[16'h021E] = 8'h00;
RAM[16'h021F] = 8'h00;
RAM[16'h0220] = 8'h00;
RAM[16'h0221] = 8'h00;
RAM[16'h0222] = 8'h00;
RAM[16'h0223] = 8'h00;
RAM[16'h0224] = 8'h00;
RAM[16'h0225] = 8'h00;
RAM[16'h0226] = 8'h00;
RAM[16'h0227] = 8'h00;
RAM[16'h0228] = 8'h00;
RAM[16'h0229] = 8'h00;
RAM[16'h022A] = 8'h00;
RAM[16'h022B] = 8'h00;
RAM[16'h022C] = 8'h00;
RAM[16'h022D] = 8'h00;
RAM[16'h022E] = 8'h00;
RAM[16'h022F] = 8'h00;
RAM[16'h0230] = 8'h00;
RAM[16'h0231] = 8'h00;
RAM[16'h0232] = 8'h00;
RAM[16'h0233] = 8'h00;
RAM[16'h0234] = 8'h00;
RAM[16'h0235] = 8'h00;
RAM[16'h0236] = 8'h00;
RAM[16'h0237] = 8'h00;
RAM[16'h0238] = 8'h00;
RAM[16'h0239] = 8'h00;
RAM[16'h023A] = 8'h00;
RAM[16'h023B] = 8'h00;
RAM[16'h023C] = 8'h00;
RAM[16'h023D] = 8'h00;
RAM[16'h023E] = 8'h00;
RAM[16'h023F] = 8'h00;
RAM[16'h0240] = 8'h00;
RAM[16'h0241] = 8'h00;
RAM[16'h0242] = 8'h00;
RAM[16'h0243] = 8'h00;
RAM[16'h0244] = 8'h00;
RAM[16'h0245] = 8'h00;
RAM[16'h0246] = 8'h00;
RAM[16'h0247] = 8'h00;
RAM[16'h0248] = 8'h00;
RAM[16'h0249] = 8'h00;
RAM[16'h024A] = 8'h00;
RAM[16'h024B] = 8'h00;
RAM[16'h024C] = 8'h00;
RAM[16'h024D] = 8'h00;
RAM[16'h024E] = 8'h00;
RAM[16'h024F] = 8'h00;
RAM[16'h0250] = 8'h00;
RAM[16'h0251] = 8'h00;
RAM[16'h0252] = 8'h00;
RAM[16'h0253] = 8'h00;
RAM[16'h0254] = 8'h00;
RAM[16'h0255] = 8'h00;
RAM[16'h0256] = 8'h00;
RAM[16'h0257] = 8'h00;
RAM[16'h0258] = 8'h00;
RAM[16'h0259] = 8'h00;
RAM[16'h025A] = 8'h00;
RAM[16'h025B] = 8'h00;
RAM[16'h025C] = 8'h00;
RAM[16'h025D] = 8'h00;
RAM[16'h025E] = 8'h00;
RAM[16'h025F] = 8'h00;
RAM[16'h0260] = 8'h00;
RAM[16'h0261] = 8'h00;
RAM[16'h0262] = 8'h00;
RAM[16'h0263] = 8'h00;
RAM[16'h0264] = 8'h00;
RAM[16'h0265] = 8'h00;
RAM[16'h0266] = 8'h00;
RAM[16'h0267] = 8'h00;
RAM[16'h0268] = 8'h00;
RAM[16'h0269] = 8'h00;
RAM[16'h026A] = 8'h00;
RAM[16'h026B] = 8'h00;
RAM[16'h026C] = 8'h00;
RAM[16'h026D] = 8'h00;
RAM[16'h026E] = 8'h00;
RAM[16'h026F] = 8'h00;
RAM[16'h0270] = 8'h00;
RAM[16'h0271] = 8'h00;
RAM[16'h0272] = 8'h00;
RAM[16'h0273] = 8'h00;
RAM[16'h0274] = 8'h00;
RAM[16'h0275] = 8'h00;
RAM[16'h0276] = 8'h00;
RAM[16'h0277] = 8'h00;
RAM[16'h0278] = 8'h00;
RAM[16'h0279] = 8'h00;
RAM[16'h027A] = 8'h00;
RAM[16'h027B] = 8'h00;
RAM[16'h027C] = 8'h00;
RAM[16'h027D] = 8'h00;
RAM[16'h027E] = 8'h00;
RAM[16'h027F] = 8'h00;
RAM[16'h0280] = 8'h00;
RAM[16'h0281] = 8'h00;
RAM[16'h0282] = 8'h00;
RAM[16'h0283] = 8'h00;
RAM[16'h0284] = 8'h00;
RAM[16'h0285] = 8'h00;
RAM[16'h0286] = 8'h00;
RAM[16'h0287] = 8'h00;
RAM[16'h0288] = 8'h00;
RAM[16'h0289] = 8'h00;
RAM[16'h028A] = 8'h00;
RAM[16'h028B] = 8'h00;
RAM[16'h028C] = 8'h00;
RAM[16'h028D] = 8'h00;
RAM[16'h028E] = 8'h00;
RAM[16'h028F] = 8'h00;
RAM[16'h0290] = 8'h00;
RAM[16'h0291] = 8'h00;
RAM[16'h0292] = 8'h00;
RAM[16'h0293] = 8'h00;
RAM[16'h0294] = 8'h00;
RAM[16'h0295] = 8'h00;
RAM[16'h0296] = 8'h00;
RAM[16'h0297] = 8'h00;
RAM[16'h0298] = 8'h00;
RAM[16'h0299] = 8'h00;
RAM[16'h029A] = 8'h00;
RAM[16'h029B] = 8'h00;
RAM[16'h029C] = 8'h00;
RAM[16'h029D] = 8'h00;
RAM[16'h029E] = 8'h00;
RAM[16'h029F] = 8'h00;
RAM[16'h02A0] = 8'h00;
RAM[16'h02A1] = 8'h00;
RAM[16'h02A2] = 8'h00;
RAM[16'h02A3] = 8'h00;
RAM[16'h02A4] = 8'h00;
RAM[16'h02A5] = 8'h00;
RAM[16'h02A6] = 8'h00;
RAM[16'h02A7] = 8'h00;
RAM[16'h02A8] = 8'h00;
RAM[16'h02A9] = 8'h00;
RAM[16'h02AA] = 8'h00;
RAM[16'h02AB] = 8'h00;
RAM[16'h02AC] = 8'h00;
RAM[16'h02AD] = 8'h00;
RAM[16'h02AE] = 8'h00;
RAM[16'h02AF] = 8'h00;
RAM[16'h02B0] = 8'h00;
RAM[16'h02B1] = 8'h00;
RAM[16'h02B2] = 8'h00;
RAM[16'h02B3] = 8'h00;
RAM[16'h02B4] = 8'h00;
RAM[16'h02B5] = 8'h00;
RAM[16'h02B6] = 8'h00;
RAM[16'h02B7] = 8'h00;
RAM[16'h02B8] = 8'h00;
RAM[16'h02B9] = 8'h00;
RAM[16'h02BA] = 8'h00;
RAM[16'h02BB] = 8'h00;
RAM[16'h02BC] = 8'h00;
RAM[16'h02BD] = 8'h00;
RAM[16'h02BE] = 8'h00;
RAM[16'h02BF] = 8'h00;
RAM[16'h02C0] = 8'h00;
RAM[16'h02C1] = 8'h00;
RAM[16'h02C2] = 8'h00;
RAM[16'h02C3] = 8'h00;
RAM[16'h02C4] = 8'h00;
RAM[16'h02C5] = 8'h00;
RAM[16'h02C6] = 8'h00;
RAM[16'h02C7] = 8'h00;
RAM[16'h02C8] = 8'h00;
RAM[16'h02C9] = 8'h00;
RAM[16'h02CA] = 8'h00;
RAM[16'h02CB] = 8'h00;
RAM[16'h02CC] = 8'h00;
RAM[16'h02CD] = 8'h00;
RAM[16'h02CE] = 8'h00;
RAM[16'h02CF] = 8'h00;
RAM[16'h02D0] = 8'h00;
RAM[16'h02D1] = 8'h00;
RAM[16'h02D2] = 8'h00;
RAM[16'h02D3] = 8'h00;
RAM[16'h02D4] = 8'h00;
RAM[16'h02D5] = 8'h00;
RAM[16'h02D6] = 8'h00;
RAM[16'h02D7] = 8'h00;
RAM[16'h02D8] = 8'h00;
RAM[16'h02D9] = 8'h00;
RAM[16'h02DA] = 8'h00;
RAM[16'h02DB] = 8'h00;
RAM[16'h02DC] = 8'h00;
RAM[16'h02DD] = 8'h00;
RAM[16'h02DE] = 8'h00;
RAM[16'h02DF] = 8'h00;
RAM[16'h02E0] = 8'h00;
RAM[16'h02E1] = 8'h00;
RAM[16'h02E2] = 8'h00;
RAM[16'h02E3] = 8'h00;
RAM[16'h02E4] = 8'h00;
RAM[16'h02E5] = 8'h00;
RAM[16'h02E6] = 8'h00;
RAM[16'h02E7] = 8'h00;
RAM[16'h02E8] = 8'h00;
RAM[16'h02E9] = 8'h00;
RAM[16'h02EA] = 8'h00;
RAM[16'h02EB] = 8'h00;
RAM[16'h02EC] = 8'h00;
RAM[16'h02ED] = 8'h00;
RAM[16'h02EE] = 8'h00;
RAM[16'h02EF] = 8'h00;
RAM[16'h02F0] = 8'h00;
RAM[16'h02F1] = 8'h00;
RAM[16'h02F2] = 8'h00;
RAM[16'h02F3] = 8'h00;
RAM[16'h02F4] = 8'h00;
RAM[16'h02F5] = 8'h00;
RAM[16'h02F6] = 8'h00;
RAM[16'h02F7] = 8'h00;
RAM[16'h02F8] = 8'h00;
RAM[16'h02F9] = 8'h00;
RAM[16'h02FA] = 8'h00;
RAM[16'h02FB] = 8'h00;
RAM[16'h02FC] = 8'h00;
RAM[16'h02FD] = 8'h00;
RAM[16'h02FE] = 8'h00;
RAM[16'h02FF] = 8'h00;
RAM[16'h0300] = 8'h00;
RAM[16'h0301] = 8'h00;
RAM[16'h0302] = 8'h00;
RAM[16'h0303] = 8'h00;
RAM[16'h0304] = 8'h00;
RAM[16'h0305] = 8'h00;
RAM[16'h0306] = 8'h00;
RAM[16'h0307] = 8'h00;
RAM[16'h0308] = 8'h00;
RAM[16'h0309] = 8'h00;
RAM[16'h030A] = 8'h00;
RAM[16'h030B] = 8'h00;
RAM[16'h030C] = 8'h00;
RAM[16'h030D] = 8'h00;
RAM[16'h030E] = 8'h00;
RAM[16'h030F] = 8'h00;
RAM[16'h0310] = 8'h00;
RAM[16'h0311] = 8'h00;
RAM[16'h0312] = 8'h00;
RAM[16'h0313] = 8'h00;
RAM[16'h0314] = 8'h00;
RAM[16'h0315] = 8'h00;
RAM[16'h0316] = 8'h00;
RAM[16'h0317] = 8'h00;
RAM[16'h0318] = 8'h00;
RAM[16'h0319] = 8'h00;
RAM[16'h031A] = 8'h00;
RAM[16'h031B] = 8'h00;
RAM[16'h031C] = 8'h00;
RAM[16'h031D] = 8'h00;
RAM[16'h031E] = 8'h00;
RAM[16'h031F] = 8'h00;
RAM[16'h0320] = 8'h00;
RAM[16'h0321] = 8'h00;
RAM[16'h0322] = 8'h00;
RAM[16'h0323] = 8'h00;
RAM[16'h0324] = 8'h00;
RAM[16'h0325] = 8'h00;
RAM[16'h0326] = 8'h00;
RAM[16'h0327] = 8'h00;
RAM[16'h0328] = 8'h00;
RAM[16'h0329] = 8'h00;
RAM[16'h032A] = 8'h00;
RAM[16'h032B] = 8'h00;
RAM[16'h032C] = 8'h00;
RAM[16'h032D] = 8'h00;
RAM[16'h032E] = 8'h00;
RAM[16'h032F] = 8'h00;
RAM[16'h0330] = 8'h00;
RAM[16'h0331] = 8'h00;
RAM[16'h0332] = 8'h00;
RAM[16'h0333] = 8'h00;
RAM[16'h0334] = 8'h00;
RAM[16'h0335] = 8'h00;
RAM[16'h0336] = 8'h00;
RAM[16'h0337] = 8'h00;
RAM[16'h0338] = 8'h00;
RAM[16'h0339] = 8'h00;
RAM[16'h033A] = 8'h00;
RAM[16'h033B] = 8'h00;
RAM[16'h033C] = 8'h00;
RAM[16'h033D] = 8'h00;
RAM[16'h033E] = 8'h00;
RAM[16'h033F] = 8'h00;
RAM[16'h0340] = 8'h00;
RAM[16'h0341] = 8'h00;
RAM[16'h0342] = 8'h00;
RAM[16'h0343] = 8'h00;
RAM[16'h0344] = 8'h00;
RAM[16'h0345] = 8'h00;
RAM[16'h0346] = 8'h00;
RAM[16'h0347] = 8'h00;
RAM[16'h0348] = 8'h00;
RAM[16'h0349] = 8'h00;
RAM[16'h034A] = 8'h00;
RAM[16'h034B] = 8'h00;
RAM[16'h034C] = 8'h00;
RAM[16'h034D] = 8'h00;
RAM[16'h034E] = 8'h00;
RAM[16'h034F] = 8'h00;
RAM[16'h0350] = 8'h00;
RAM[16'h0351] = 8'h00;
RAM[16'h0352] = 8'h00;
RAM[16'h0353] = 8'h00;
RAM[16'h0354] = 8'h00;
RAM[16'h0355] = 8'h00;
RAM[16'h0356] = 8'h00;
RAM[16'h0357] = 8'h00;
RAM[16'h0358] = 8'h00;
RAM[16'h0359] = 8'h00;
RAM[16'h035A] = 8'h00;
RAM[16'h035B] = 8'h00;
RAM[16'h035C] = 8'h00;
RAM[16'h035D] = 8'h00;
RAM[16'h035E] = 8'h00;
RAM[16'h035F] = 8'h00;
RAM[16'h0360] = 8'h00;
RAM[16'h0361] = 8'h00;
RAM[16'h0362] = 8'h00;
RAM[16'h0363] = 8'h00;
RAM[16'h0364] = 8'h00;
RAM[16'h0365] = 8'h00;
RAM[16'h0366] = 8'h00;
RAM[16'h0367] = 8'h00;
RAM[16'h0368] = 8'h00;
RAM[16'h0369] = 8'h00;
RAM[16'h036A] = 8'h00;
RAM[16'h036B] = 8'h00;
RAM[16'h036C] = 8'h00;
RAM[16'h036D] = 8'h00;
RAM[16'h036E] = 8'h00;
RAM[16'h036F] = 8'h00;
RAM[16'h0370] = 8'h00;
RAM[16'h0371] = 8'h00;
RAM[16'h0372] = 8'h00;
RAM[16'h0373] = 8'h00;
RAM[16'h0374] = 8'h00;
RAM[16'h0375] = 8'h00;
RAM[16'h0376] = 8'h00;
RAM[16'h0377] = 8'h00;
RAM[16'h0378] = 8'h00;
RAM[16'h0379] = 8'h00;
RAM[16'h037A] = 8'h00;
RAM[16'h037B] = 8'h00;
RAM[16'h037C] = 8'h00;
RAM[16'h037D] = 8'h00;
RAM[16'h037E] = 8'h00;
RAM[16'h037F] = 8'h00;
RAM[16'h0380] = 8'h00;
RAM[16'h0381] = 8'h00;
RAM[16'h0382] = 8'h00;
RAM[16'h0383] = 8'h00;
RAM[16'h0384] = 8'h00;
RAM[16'h0385] = 8'h00;
RAM[16'h0386] = 8'h00;
RAM[16'h0387] = 8'h00;
RAM[16'h0388] = 8'h00;
RAM[16'h0389] = 8'h00;
RAM[16'h038A] = 8'h00;
RAM[16'h038B] = 8'h00;
RAM[16'h038C] = 8'h00;
RAM[16'h038D] = 8'h00;
RAM[16'h038E] = 8'h00;
RAM[16'h038F] = 8'h00;
RAM[16'h0390] = 8'h00;
RAM[16'h0391] = 8'h00;
RAM[16'h0392] = 8'h00;
RAM[16'h0393] = 8'h00;
RAM[16'h0394] = 8'h00;
RAM[16'h0395] = 8'h00;
RAM[16'h0396] = 8'h00;
RAM[16'h0397] = 8'h00;
RAM[16'h0398] = 8'h00;
RAM[16'h0399] = 8'h00;
RAM[16'h039A] = 8'h00;
RAM[16'h039B] = 8'h00;
RAM[16'h039C] = 8'h00;
RAM[16'h039D] = 8'h00;
RAM[16'h039E] = 8'h00;
RAM[16'h039F] = 8'h00;
RAM[16'h03A0] = 8'h00;
RAM[16'h03A1] = 8'h00;
RAM[16'h03A2] = 8'h00;
RAM[16'h03A3] = 8'h00;
RAM[16'h03A4] = 8'h00;
RAM[16'h03A5] = 8'h00;
RAM[16'h03A6] = 8'h00;
RAM[16'h03A7] = 8'h00;
RAM[16'h03A8] = 8'h00;
RAM[16'h03A9] = 8'h00;
RAM[16'h03AA] = 8'h00;
RAM[16'h03AB] = 8'h00;
RAM[16'h03AC] = 8'h00;
RAM[16'h03AD] = 8'h00;
RAM[16'h03AE] = 8'h00;
RAM[16'h03AF] = 8'h00;
RAM[16'h03B0] = 8'h00;
RAM[16'h03B1] = 8'h00;
RAM[16'h03B2] = 8'h00;
RAM[16'h03B3] = 8'h00;
RAM[16'h03B4] = 8'h00;
RAM[16'h03B5] = 8'h00;
RAM[16'h03B6] = 8'h00;
RAM[16'h03B7] = 8'h00;
RAM[16'h03B8] = 8'h00;
RAM[16'h03B9] = 8'h00;
RAM[16'h03BA] = 8'h00;
RAM[16'h03BB] = 8'h00;
RAM[16'h03BC] = 8'h00;
RAM[16'h03BD] = 8'h00;
RAM[16'h03BE] = 8'h00;
RAM[16'h03BF] = 8'h00;
RAM[16'h03C0] = 8'h00;
RAM[16'h03C1] = 8'h00;
RAM[16'h03C2] = 8'h00;
RAM[16'h03C3] = 8'h00;
RAM[16'h03C4] = 8'h00;
RAM[16'h03C5] = 8'h00;
RAM[16'h03C6] = 8'h00;
RAM[16'h03C7] = 8'h00;
RAM[16'h03C8] = 8'h00;
RAM[16'h03C9] = 8'h00;
RAM[16'h03CA] = 8'h00;
RAM[16'h03CB] = 8'h00;
RAM[16'h03CC] = 8'h00;
RAM[16'h03CD] = 8'h00;
RAM[16'h03CE] = 8'h00;
RAM[16'h03CF] = 8'h00;
RAM[16'h03D0] = 8'h00;
RAM[16'h03D1] = 8'h00;
RAM[16'h03D2] = 8'h00;
RAM[16'h03D3] = 8'h00;
RAM[16'h03D4] = 8'h00;
RAM[16'h03D5] = 8'h00;
RAM[16'h03D6] = 8'h00;
RAM[16'h03D7] = 8'h00;
RAM[16'h03D8] = 8'h00;
RAM[16'h03D9] = 8'h00;
RAM[16'h03DA] = 8'h00;
RAM[16'h03DB] = 8'h00;
RAM[16'h03DC] = 8'h00;
RAM[16'h03DD] = 8'h00;
RAM[16'h03DE] = 8'h00;
RAM[16'h03DF] = 8'h00;
RAM[16'h03E0] = 8'h00;
RAM[16'h03E1] = 8'h00;
RAM[16'h03E2] = 8'h00;
RAM[16'h03E3] = 8'h00;
RAM[16'h03E4] = 8'h00;
RAM[16'h03E5] = 8'h00;
RAM[16'h03E6] = 8'h00;
RAM[16'h03E7] = 8'h00;
RAM[16'h03E8] = 8'h00;
RAM[16'h03E9] = 8'h00;
RAM[16'h03EA] = 8'h00;
RAM[16'h03EB] = 8'h00;
RAM[16'h03EC] = 8'h00;
RAM[16'h03ED] = 8'h00;
RAM[16'h03EE] = 8'h00;
RAM[16'h03EF] = 8'h00;
RAM[16'h03F0] = 8'h00;
RAM[16'h03F1] = 8'h00;
RAM[16'h03F2] = 8'h00;
RAM[16'h03F3] = 8'h00;
RAM[16'h03F4] = 8'h00;
RAM[16'h03F5] = 8'h00;
RAM[16'h03F6] = 8'h00;
RAM[16'h03F7] = 8'h00;
RAM[16'h03F8] = 8'h00;
RAM[16'h03F9] = 8'h00;
RAM[16'h03FA] = 8'h00;
RAM[16'h03FB] = 8'h00;
RAM[16'h03FC] = 8'h00;
RAM[16'h03FD] = 8'h00;
RAM[16'h03FE] = 8'h00;
RAM[16'h03FF] = 8'h00;
RAM[16'h0400] = 8'h00;
RAM[16'h0401] = 8'h00;
RAM[16'h0402] = 8'h00;
RAM[16'h0403] = 8'h00;
RAM[16'h0404] = 8'h00;
RAM[16'h0405] = 8'h00;
RAM[16'h0406] = 8'h00;
RAM[16'h0407] = 8'h00;
RAM[16'h0408] = 8'h00;
RAM[16'h0409] = 8'h00;
RAM[16'h040A] = 8'h00;
RAM[16'h040B] = 8'h00;
RAM[16'h040C] = 8'h00;
RAM[16'h040D] = 8'h00;
RAM[16'h040E] = 8'h00;
RAM[16'h040F] = 8'h00;
RAM[16'h0410] = 8'h00;
RAM[16'h0411] = 8'h00;
RAM[16'h0412] = 8'h00;
RAM[16'h0413] = 8'h00;
RAM[16'h0414] = 8'h00;
RAM[16'h0415] = 8'h00;
RAM[16'h0416] = 8'h00;
RAM[16'h0417] = 8'h00;
RAM[16'h0418] = 8'h00;
RAM[16'h0419] = 8'h00;
RAM[16'h041A] = 8'h00;
RAM[16'h041B] = 8'h00;
RAM[16'h041C] = 8'h00;
RAM[16'h041D] = 8'h00;
RAM[16'h041E] = 8'h00;
RAM[16'h041F] = 8'h00;
RAM[16'h0420] = 8'h00;
RAM[16'h0421] = 8'h00;
RAM[16'h0422] = 8'h00;
RAM[16'h0423] = 8'h00;
RAM[16'h0424] = 8'h00;
RAM[16'h0425] = 8'h00;
RAM[16'h0426] = 8'h00;
RAM[16'h0427] = 8'h00;
RAM[16'h0428] = 8'h00;
RAM[16'h0429] = 8'h00;
RAM[16'h042A] = 8'h00;
RAM[16'h042B] = 8'h00;
RAM[16'h042C] = 8'h00;
RAM[16'h042D] = 8'h00;
RAM[16'h042E] = 8'h00;
RAM[16'h042F] = 8'h00;
RAM[16'h0430] = 8'h00;
RAM[16'h0431] = 8'h00;
RAM[16'h0432] = 8'h00;
RAM[16'h0433] = 8'h00;
RAM[16'h0434] = 8'h00;
RAM[16'h0435] = 8'h00;
RAM[16'h0436] = 8'h00;
RAM[16'h0437] = 8'h00;
RAM[16'h0438] = 8'h00;
RAM[16'h0439] = 8'h00;
RAM[16'h043A] = 8'h00;
RAM[16'h043B] = 8'h00;
RAM[16'h043C] = 8'h00;
RAM[16'h043D] = 8'h00;
RAM[16'h043E] = 8'h00;
RAM[16'h043F] = 8'h00;
RAM[16'h0440] = 8'h00;
RAM[16'h0441] = 8'h00;
RAM[16'h0442] = 8'h00;
RAM[16'h0443] = 8'h00;
RAM[16'h0444] = 8'h00;
RAM[16'h0445] = 8'h00;
RAM[16'h0446] = 8'h00;
RAM[16'h0447] = 8'h00;
RAM[16'h0448] = 8'h00;
RAM[16'h0449] = 8'h00;
RAM[16'h044A] = 8'h00;
RAM[16'h044B] = 8'h00;
RAM[16'h044C] = 8'h00;
RAM[16'h044D] = 8'h00;
RAM[16'h044E] = 8'h00;
RAM[16'h044F] = 8'h00;
RAM[16'h0450] = 8'h00;
RAM[16'h0451] = 8'h00;
RAM[16'h0452] = 8'h00;
RAM[16'h0453] = 8'h00;
RAM[16'h0454] = 8'h00;
RAM[16'h0455] = 8'h00;
RAM[16'h0456] = 8'h00;
RAM[16'h0457] = 8'h00;
RAM[16'h0458] = 8'h00;
RAM[16'h0459] = 8'h00;
RAM[16'h045A] = 8'h00;
RAM[16'h045B] = 8'h00;
RAM[16'h045C] = 8'h00;
RAM[16'h045D] = 8'h00;
RAM[16'h045E] = 8'h00;
RAM[16'h045F] = 8'h00;
RAM[16'h0460] = 8'h00;
RAM[16'h0461] = 8'h00;
RAM[16'h0462] = 8'h00;
RAM[16'h0463] = 8'h00;
RAM[16'h0464] = 8'h00;
RAM[16'h0465] = 8'h00;
RAM[16'h0466] = 8'h00;
RAM[16'h0467] = 8'h00;
RAM[16'h0468] = 8'h00;
RAM[16'h0469] = 8'h00;
RAM[16'h046A] = 8'h00;
RAM[16'h046B] = 8'h00;
RAM[16'h046C] = 8'h00;
RAM[16'h046D] = 8'h00;
RAM[16'h046E] = 8'h00;
RAM[16'h046F] = 8'h00;
RAM[16'h0470] = 8'h00;
RAM[16'h0471] = 8'h00;
RAM[16'h0472] = 8'h00;
RAM[16'h0473] = 8'h00;
RAM[16'h0474] = 8'h00;
RAM[16'h0475] = 8'h00;
RAM[16'h0476] = 8'h00;
RAM[16'h0477] = 8'h00;
RAM[16'h0478] = 8'h00;
RAM[16'h0479] = 8'h00;
RAM[16'h047A] = 8'h00;
RAM[16'h047B] = 8'h00;
RAM[16'h047C] = 8'h00;
RAM[16'h047D] = 8'h00;
RAM[16'h047E] = 8'h00;
RAM[16'h047F] = 8'h00;
RAM[16'h0480] = 8'h00;
RAM[16'h0481] = 8'h00;
RAM[16'h0482] = 8'h00;
RAM[16'h0483] = 8'h00;
RAM[16'h0484] = 8'h00;
RAM[16'h0485] = 8'h00;
RAM[16'h0486] = 8'h00;
RAM[16'h0487] = 8'h00;
RAM[16'h0488] = 8'h00;
RAM[16'h0489] = 8'h00;
RAM[16'h048A] = 8'h00;
RAM[16'h048B] = 8'h00;
RAM[16'h048C] = 8'h00;
RAM[16'h048D] = 8'h00;
RAM[16'h048E] = 8'h00;
RAM[16'h048F] = 8'h00;
RAM[16'h0490] = 8'h00;
RAM[16'h0491] = 8'h00;
RAM[16'h0492] = 8'h00;
RAM[16'h0493] = 8'h00;
RAM[16'h0494] = 8'h00;
RAM[16'h0495] = 8'h00;
RAM[16'h0496] = 8'h00;
RAM[16'h0497] = 8'h00;
RAM[16'h0498] = 8'h00;
RAM[16'h0499] = 8'h00;
RAM[16'h049A] = 8'h00;
RAM[16'h049B] = 8'h00;
RAM[16'h049C] = 8'h00;
RAM[16'h049D] = 8'h00;
RAM[16'h049E] = 8'h00;
RAM[16'h049F] = 8'h00;
RAM[16'h04A0] = 8'h00;
RAM[16'h04A1] = 8'h00;
RAM[16'h04A2] = 8'h00;
RAM[16'h04A3] = 8'h00;
RAM[16'h04A4] = 8'h00;
RAM[16'h04A5] = 8'h00;
RAM[16'h04A6] = 8'h00;
RAM[16'h04A7] = 8'h00;
RAM[16'h04A8] = 8'h00;
RAM[16'h04A9] = 8'h00;
RAM[16'h04AA] = 8'h00;
RAM[16'h04AB] = 8'h00;
RAM[16'h04AC] = 8'h00;
RAM[16'h04AD] = 8'h00;
RAM[16'h04AE] = 8'h00;
RAM[16'h04AF] = 8'h00;
RAM[16'h04B0] = 8'h00;
RAM[16'h04B1] = 8'h00;
RAM[16'h04B2] = 8'h00;
RAM[16'h04B3] = 8'h00;
RAM[16'h04B4] = 8'h00;
RAM[16'h04B5] = 8'h00;
RAM[16'h04B6] = 8'h00;
RAM[16'h04B7] = 8'h00;
RAM[16'h04B8] = 8'h00;
RAM[16'h04B9] = 8'h00;
RAM[16'h04BA] = 8'h00;
RAM[16'h04BB] = 8'h00;
RAM[16'h04BC] = 8'h00;
RAM[16'h04BD] = 8'h00;
RAM[16'h04BE] = 8'h00;
RAM[16'h04BF] = 8'h00;
RAM[16'h04C0] = 8'h00;
RAM[16'h04C1] = 8'h00;
RAM[16'h04C2] = 8'h00;
RAM[16'h04C3] = 8'h00;
RAM[16'h04C4] = 8'h00;
RAM[16'h04C5] = 8'h00;
RAM[16'h04C6] = 8'h00;
RAM[16'h04C7] = 8'h00;
RAM[16'h04C8] = 8'h00;
RAM[16'h04C9] = 8'h00;
RAM[16'h04CA] = 8'h00;
RAM[16'h04CB] = 8'h00;
RAM[16'h04CC] = 8'h00;
RAM[16'h04CD] = 8'h00;
RAM[16'h04CE] = 8'h00;
RAM[16'h04CF] = 8'h00;
RAM[16'h04D0] = 8'h00;
RAM[16'h04D1] = 8'h00;
RAM[16'h04D2] = 8'h00;
RAM[16'h04D3] = 8'h00;
RAM[16'h04D4] = 8'h00;
RAM[16'h04D5] = 8'h00;
RAM[16'h04D6] = 8'h00;
RAM[16'h04D7] = 8'h00;
RAM[16'h04D8] = 8'h00;
RAM[16'h04D9] = 8'h00;
RAM[16'h04DA] = 8'h00;
RAM[16'h04DB] = 8'h00;
RAM[16'h04DC] = 8'h00;
RAM[16'h04DD] = 8'h00;
RAM[16'h04DE] = 8'h00;
RAM[16'h04DF] = 8'h00;
RAM[16'h04E0] = 8'h00;
RAM[16'h04E1] = 8'h00;
RAM[16'h04E2] = 8'h00;
RAM[16'h04E3] = 8'h00;
RAM[16'h04E4] = 8'h00;
RAM[16'h04E5] = 8'h00;
RAM[16'h04E6] = 8'h00;
RAM[16'h04E7] = 8'h00;
RAM[16'h04E8] = 8'h00;
RAM[16'h04E9] = 8'h00;
RAM[16'h04EA] = 8'h00;
RAM[16'h04EB] = 8'h00;
RAM[16'h04EC] = 8'h00;
RAM[16'h04ED] = 8'h00;
RAM[16'h04EE] = 8'h00;
RAM[16'h04EF] = 8'h00;
RAM[16'h04F0] = 8'h00;
RAM[16'h04F1] = 8'h00;
RAM[16'h04F2] = 8'h00;
RAM[16'h04F3] = 8'h00;
RAM[16'h04F4] = 8'h00;
RAM[16'h04F5] = 8'h00;
RAM[16'h04F6] = 8'h00;
RAM[16'h04F7] = 8'h00;
RAM[16'h04F8] = 8'h00;
RAM[16'h04F9] = 8'h00;
RAM[16'h04FA] = 8'h00;
RAM[16'h04FB] = 8'h00;
RAM[16'h04FC] = 8'h00;
RAM[16'h04FD] = 8'h00;
RAM[16'h04FE] = 8'h00;
RAM[16'h04FF] = 8'h00;
RAM[16'h0500] = 8'h00;
RAM[16'h0501] = 8'h00;
RAM[16'h0502] = 8'h00;
RAM[16'h0503] = 8'h00;
RAM[16'h0504] = 8'h00;
RAM[16'h0505] = 8'h00;
RAM[16'h0506] = 8'h00;
RAM[16'h0507] = 8'h00;
RAM[16'h0508] = 8'h00;
RAM[16'h0509] = 8'h00;
RAM[16'h050A] = 8'h00;
RAM[16'h050B] = 8'h00;
RAM[16'h050C] = 8'h00;
RAM[16'h050D] = 8'h00;
RAM[16'h050E] = 8'h00;
RAM[16'h050F] = 8'h00;
RAM[16'h0510] = 8'h00;
RAM[16'h0511] = 8'h00;
RAM[16'h0512] = 8'h00;
RAM[16'h0513] = 8'h00;
RAM[16'h0514] = 8'h00;
RAM[16'h0515] = 8'h00;
RAM[16'h0516] = 8'h00;
RAM[16'h0517] = 8'h00;
RAM[16'h0518] = 8'h00;
RAM[16'h0519] = 8'h00;
RAM[16'h051A] = 8'h00;
RAM[16'h051B] = 8'h00;
RAM[16'h051C] = 8'h00;
RAM[16'h051D] = 8'h00;
RAM[16'h051E] = 8'h00;
RAM[16'h051F] = 8'h00;
RAM[16'h0520] = 8'h00;
RAM[16'h0521] = 8'h00;
RAM[16'h0522] = 8'h00;
RAM[16'h0523] = 8'h00;
RAM[16'h0524] = 8'h00;
RAM[16'h0525] = 8'h00;
RAM[16'h0526] = 8'h00;
RAM[16'h0527] = 8'h00;
RAM[16'h0528] = 8'h00;
RAM[16'h0529] = 8'h00;
RAM[16'h052A] = 8'h00;
RAM[16'h052B] = 8'h00;
RAM[16'h052C] = 8'h00;
RAM[16'h052D] = 8'h00;
RAM[16'h052E] = 8'h00;
RAM[16'h052F] = 8'h00;
RAM[16'h0530] = 8'h00;
RAM[16'h0531] = 8'h00;
RAM[16'h0532] = 8'h00;
RAM[16'h0533] = 8'h00;
RAM[16'h0534] = 8'h00;
RAM[16'h0535] = 8'h00;
RAM[16'h0536] = 8'h00;
RAM[16'h0537] = 8'h00;
RAM[16'h0538] = 8'h00;
RAM[16'h0539] = 8'h00;
RAM[16'h053A] = 8'h00;
RAM[16'h053B] = 8'h00;
RAM[16'h053C] = 8'h00;
RAM[16'h053D] = 8'h00;
RAM[16'h053E] = 8'h00;
RAM[16'h053F] = 8'h00;
RAM[16'h0540] = 8'h00;
RAM[16'h0541] = 8'h00;
RAM[16'h0542] = 8'h00;
RAM[16'h0543] = 8'h00;
RAM[16'h0544] = 8'h00;
RAM[16'h0545] = 8'h00;
RAM[16'h0546] = 8'h00;
RAM[16'h0547] = 8'h00;
RAM[16'h0548] = 8'h00;
RAM[16'h0549] = 8'h00;
RAM[16'h054A] = 8'h00;
RAM[16'h054B] = 8'h00;
RAM[16'h054C] = 8'h00;
RAM[16'h054D] = 8'h00;
RAM[16'h054E] = 8'h00;
RAM[16'h054F] = 8'h00;
RAM[16'h0550] = 8'h00;
RAM[16'h0551] = 8'h00;
RAM[16'h0552] = 8'h00;
RAM[16'h0553] = 8'h00;
RAM[16'h0554] = 8'h00;
RAM[16'h0555] = 8'h00;
RAM[16'h0556] = 8'h00;
RAM[16'h0557] = 8'h00;
RAM[16'h0558] = 8'h00;
RAM[16'h0559] = 8'h00;
RAM[16'h055A] = 8'h00;
RAM[16'h055B] = 8'h00;
RAM[16'h055C] = 8'h00;
RAM[16'h055D] = 8'h00;
RAM[16'h055E] = 8'h00;
RAM[16'h055F] = 8'h00;
RAM[16'h0560] = 8'h00;
RAM[16'h0561] = 8'h00;
RAM[16'h0562] = 8'h00;
RAM[16'h0563] = 8'h00;
RAM[16'h0564] = 8'h00;
RAM[16'h0565] = 8'h00;
RAM[16'h0566] = 8'h00;
RAM[16'h0567] = 8'h00;
RAM[16'h0568] = 8'h00;
RAM[16'h0569] = 8'h00;
RAM[16'h056A] = 8'h00;
RAM[16'h056B] = 8'h00;
RAM[16'h056C] = 8'h00;
RAM[16'h056D] = 8'h00;
RAM[16'h056E] = 8'h00;
RAM[16'h056F] = 8'h00;
RAM[16'h0570] = 8'h00;
RAM[16'h0571] = 8'h00;
RAM[16'h0572] = 8'h00;
RAM[16'h0573] = 8'h00;
RAM[16'h0574] = 8'h00;
RAM[16'h0575] = 8'h00;
RAM[16'h0576] = 8'h00;
RAM[16'h0577] = 8'h00;
RAM[16'h0578] = 8'h00;
RAM[16'h0579] = 8'h00;
RAM[16'h057A] = 8'h00;
RAM[16'h057B] = 8'h00;
RAM[16'h057C] = 8'h00;
RAM[16'h057D] = 8'h00;
RAM[16'h057E] = 8'h00;
RAM[16'h057F] = 8'h00;
RAM[16'h0580] = 8'h00;
RAM[16'h0581] = 8'h00;
RAM[16'h0582] = 8'h00;
RAM[16'h0583] = 8'h00;
RAM[16'h0584] = 8'h00;
RAM[16'h0585] = 8'h00;
RAM[16'h0586] = 8'h00;
RAM[16'h0587] = 8'h00;
RAM[16'h0588] = 8'h00;
RAM[16'h0589] = 8'h00;
RAM[16'h058A] = 8'h00;
RAM[16'h058B] = 8'h00;
RAM[16'h058C] = 8'h00;
RAM[16'h058D] = 8'h00;
RAM[16'h058E] = 8'h00;
RAM[16'h058F] = 8'h00;
RAM[16'h0590] = 8'h00;
RAM[16'h0591] = 8'h00;
RAM[16'h0592] = 8'h00;
RAM[16'h0593] = 8'h00;
RAM[16'h0594] = 8'h00;
RAM[16'h0595] = 8'h00;
RAM[16'h0596] = 8'h00;
RAM[16'h0597] = 8'h00;
RAM[16'h0598] = 8'h00;
RAM[16'h0599] = 8'h00;
RAM[16'h059A] = 8'h00;
RAM[16'h059B] = 8'h00;
RAM[16'h059C] = 8'h00;
RAM[16'h059D] = 8'h00;
RAM[16'h059E] = 8'h00;
RAM[16'h059F] = 8'h00;
RAM[16'h05A0] = 8'h00;
RAM[16'h05A1] = 8'h00;
RAM[16'h05A2] = 8'h00;
RAM[16'h05A3] = 8'h00;
RAM[16'h05A4] = 8'h00;
RAM[16'h05A5] = 8'h00;
RAM[16'h05A6] = 8'h00;
RAM[16'h05A7] = 8'h00;
RAM[16'h05A8] = 8'h00;
RAM[16'h05A9] = 8'h00;
RAM[16'h05AA] = 8'h00;
RAM[16'h05AB] = 8'h00;
RAM[16'h05AC] = 8'h00;
RAM[16'h05AD] = 8'h00;
RAM[16'h05AE] = 8'h00;
RAM[16'h05AF] = 8'h00;
RAM[16'h05B0] = 8'h00;
RAM[16'h05B1] = 8'h00;
RAM[16'h05B2] = 8'h00;
RAM[16'h05B3] = 8'h00;
RAM[16'h05B4] = 8'h00;
RAM[16'h05B5] = 8'h00;
RAM[16'h05B6] = 8'h00;
RAM[16'h05B7] = 8'h00;
RAM[16'h05B8] = 8'h00;
RAM[16'h05B9] = 8'h00;
RAM[16'h05BA] = 8'h00;
RAM[16'h05BB] = 8'h00;
RAM[16'h05BC] = 8'h00;
RAM[16'h05BD] = 8'h00;
RAM[16'h05BE] = 8'h00;
RAM[16'h05BF] = 8'h00;
RAM[16'h05C0] = 8'h00;
RAM[16'h05C1] = 8'h00;
RAM[16'h05C2] = 8'h00;
RAM[16'h05C3] = 8'h00;
RAM[16'h05C4] = 8'h00;
RAM[16'h05C5] = 8'h00;
RAM[16'h05C6] = 8'h00;
RAM[16'h05C7] = 8'h00;
RAM[16'h05C8] = 8'h00;
RAM[16'h05C9] = 8'h00;
RAM[16'h05CA] = 8'h00;
RAM[16'h05CB] = 8'h00;
RAM[16'h05CC] = 8'h00;
RAM[16'h05CD] = 8'h00;
RAM[16'h05CE] = 8'h00;
RAM[16'h05CF] = 8'h00;
RAM[16'h05D0] = 8'h00;
RAM[16'h05D1] = 8'h00;
RAM[16'h05D2] = 8'h00;
RAM[16'h05D3] = 8'h00;
RAM[16'h05D4] = 8'h00;
RAM[16'h05D5] = 8'h00;
RAM[16'h05D6] = 8'h00;
RAM[16'h05D7] = 8'h00;
RAM[16'h05D8] = 8'h00;
RAM[16'h05D9] = 8'h00;
RAM[16'h05DA] = 8'h00;
RAM[16'h05DB] = 8'h00;
RAM[16'h05DC] = 8'h00;
RAM[16'h05DD] = 8'h00;
RAM[16'h05DE] = 8'h00;
RAM[16'h05DF] = 8'h00;
RAM[16'h05E0] = 8'h00;
RAM[16'h05E1] = 8'h00;
RAM[16'h05E2] = 8'h00;
RAM[16'h05E3] = 8'h00;
RAM[16'h05E4] = 8'h00;
RAM[16'h05E5] = 8'h00;
RAM[16'h05E6] = 8'h00;
RAM[16'h05E7] = 8'h00;
RAM[16'h05E8] = 8'h00;
RAM[16'h05E9] = 8'h00;
RAM[16'h05EA] = 8'h00;
RAM[16'h05EB] = 8'h00;
RAM[16'h05EC] = 8'h00;
RAM[16'h05ED] = 8'h00;
RAM[16'h05EE] = 8'h00;
RAM[16'h05EF] = 8'h00;
RAM[16'h05F0] = 8'h00;
RAM[16'h05F1] = 8'h00;
RAM[16'h05F2] = 8'h00;
RAM[16'h05F3] = 8'h00;
RAM[16'h05F4] = 8'h00;
RAM[16'h05F5] = 8'h00;
RAM[16'h05F6] = 8'h00;
RAM[16'h05F7] = 8'h00;
RAM[16'h05F8] = 8'h00;
RAM[16'h05F9] = 8'h00;
RAM[16'h05FA] = 8'h00;
RAM[16'h05FB] = 8'h00;
RAM[16'h05FC] = 8'h00;
RAM[16'h05FD] = 8'h00;
RAM[16'h05FE] = 8'h00;
RAM[16'h05FF] = 8'h00;
RAM[16'h0600] = 8'h00;
RAM[16'h0601] = 8'h00;
RAM[16'h0602] = 8'h00;
RAM[16'h0603] = 8'h00;
RAM[16'h0604] = 8'h00;
RAM[16'h0605] = 8'h00;
RAM[16'h0606] = 8'h00;
RAM[16'h0607] = 8'h00;
RAM[16'h0608] = 8'h00;
RAM[16'h0609] = 8'h00;
RAM[16'h060A] = 8'h00;
RAM[16'h060B] = 8'h00;
RAM[16'h060C] = 8'h00;
RAM[16'h060D] = 8'h00;
RAM[16'h060E] = 8'h00;
RAM[16'h060F] = 8'h00;
RAM[16'h0610] = 8'h00;
RAM[16'h0611] = 8'h00;
RAM[16'h0612] = 8'h00;
RAM[16'h0613] = 8'h00;
RAM[16'h0614] = 8'h00;
RAM[16'h0615] = 8'h00;
RAM[16'h0616] = 8'h00;
RAM[16'h0617] = 8'h00;
RAM[16'h0618] = 8'h00;
RAM[16'h0619] = 8'h00;
RAM[16'h061A] = 8'h00;
RAM[16'h061B] = 8'h00;
RAM[16'h061C] = 8'h00;
RAM[16'h061D] = 8'h00;
RAM[16'h061E] = 8'h00;
RAM[16'h061F] = 8'h00;
RAM[16'h0620] = 8'h00;
RAM[16'h0621] = 8'h00;
RAM[16'h0622] = 8'h00;
RAM[16'h0623] = 8'h00;
RAM[16'h0624] = 8'h00;
RAM[16'h0625] = 8'h00;
RAM[16'h0626] = 8'h00;
RAM[16'h0627] = 8'h00;
RAM[16'h0628] = 8'h00;
RAM[16'h0629] = 8'h00;
RAM[16'h062A] = 8'h00;
RAM[16'h062B] = 8'h00;
RAM[16'h062C] = 8'h00;
RAM[16'h062D] = 8'h00;
RAM[16'h062E] = 8'h00;
RAM[16'h062F] = 8'h00;
RAM[16'h0630] = 8'h00;
RAM[16'h0631] = 8'h00;
RAM[16'h0632] = 8'h00;
RAM[16'h0633] = 8'h00;
RAM[16'h0634] = 8'h00;
RAM[16'h0635] = 8'h00;
RAM[16'h0636] = 8'h00;
RAM[16'h0637] = 8'h00;
RAM[16'h0638] = 8'h00;
RAM[16'h0639] = 8'h00;
RAM[16'h063A] = 8'h00;
RAM[16'h063B] = 8'h00;
RAM[16'h063C] = 8'h00;
RAM[16'h063D] = 8'h00;
RAM[16'h063E] = 8'h00;
RAM[16'h063F] = 8'h00;
RAM[16'h0640] = 8'h00;
RAM[16'h0641] = 8'h00;
RAM[16'h0642] = 8'h00;
RAM[16'h0643] = 8'h00;
RAM[16'h0644] = 8'h00;
RAM[16'h0645] = 8'h00;
RAM[16'h0646] = 8'h00;
RAM[16'h0647] = 8'h00;
RAM[16'h0648] = 8'h00;
RAM[16'h0649] = 8'h00;
RAM[16'h064A] = 8'h00;
RAM[16'h064B] = 8'h00;
RAM[16'h064C] = 8'h00;
RAM[16'h064D] = 8'h00;
RAM[16'h064E] = 8'h00;
RAM[16'h064F] = 8'h00;
RAM[16'h0650] = 8'h00;
RAM[16'h0651] = 8'h00;
RAM[16'h0652] = 8'h00;
RAM[16'h0653] = 8'h00;
RAM[16'h0654] = 8'h00;
RAM[16'h0655] = 8'h00;
RAM[16'h0656] = 8'h00;
RAM[16'h0657] = 8'h00;
RAM[16'h0658] = 8'h00;
RAM[16'h0659] = 8'h00;
RAM[16'h065A] = 8'h00;
RAM[16'h065B] = 8'h00;
RAM[16'h065C] = 8'h00;
RAM[16'h065D] = 8'h00;
RAM[16'h065E] = 8'h00;
RAM[16'h065F] = 8'h00;
RAM[16'h0660] = 8'h00;
RAM[16'h0661] = 8'h00;
RAM[16'h0662] = 8'h00;
RAM[16'h0663] = 8'h00;
RAM[16'h0664] = 8'h00;
RAM[16'h0665] = 8'h00;
RAM[16'h0666] = 8'h00;
RAM[16'h0667] = 8'h00;
RAM[16'h0668] = 8'h00;
RAM[16'h0669] = 8'h00;
RAM[16'h066A] = 8'h00;
RAM[16'h066B] = 8'h00;
RAM[16'h066C] = 8'h00;
RAM[16'h066D] = 8'h00;
RAM[16'h066E] = 8'h00;
RAM[16'h066F] = 8'h00;
RAM[16'h0670] = 8'h00;
RAM[16'h0671] = 8'h00;
RAM[16'h0672] = 8'h00;
RAM[16'h0673] = 8'h00;
RAM[16'h0674] = 8'h00;
RAM[16'h0675] = 8'h00;
RAM[16'h0676] = 8'h00;
RAM[16'h0677] = 8'h00;
RAM[16'h0678] = 8'h00;
RAM[16'h0679] = 8'h00;
RAM[16'h067A] = 8'h00;
RAM[16'h067B] = 8'h00;
RAM[16'h067C] = 8'h00;
RAM[16'h067D] = 8'h00;
RAM[16'h067E] = 8'h00;
RAM[16'h067F] = 8'h00;
RAM[16'h0680] = 8'h00;
RAM[16'h0681] = 8'h00;
RAM[16'h0682] = 8'h00;
RAM[16'h0683] = 8'h00;
RAM[16'h0684] = 8'h00;
RAM[16'h0685] = 8'h00;
RAM[16'h0686] = 8'h00;
RAM[16'h0687] = 8'h00;
RAM[16'h0688] = 8'h00;
RAM[16'h0689] = 8'h00;
RAM[16'h068A] = 8'h00;
RAM[16'h068B] = 8'h00;
RAM[16'h068C] = 8'h00;
RAM[16'h068D] = 8'h00;
RAM[16'h068E] = 8'h00;
RAM[16'h068F] = 8'h00;
RAM[16'h0690] = 8'h00;
RAM[16'h0691] = 8'h00;
RAM[16'h0692] = 8'h00;
RAM[16'h0693] = 8'h00;
RAM[16'h0694] = 8'h00;
RAM[16'h0695] = 8'h00;
RAM[16'h0696] = 8'h00;
RAM[16'h0697] = 8'h00;
RAM[16'h0698] = 8'h00;
RAM[16'h0699] = 8'h00;
RAM[16'h069A] = 8'h00;
RAM[16'h069B] = 8'h00;
RAM[16'h069C] = 8'h00;
RAM[16'h069D] = 8'h00;
RAM[16'h069E] = 8'h00;
RAM[16'h069F] = 8'h00;
RAM[16'h06A0] = 8'h00;
RAM[16'h06A1] = 8'h00;
RAM[16'h06A2] = 8'h00;
RAM[16'h06A3] = 8'h00;
RAM[16'h06A4] = 8'h00;
RAM[16'h06A5] = 8'h00;
RAM[16'h06A6] = 8'h00;
RAM[16'h06A7] = 8'h00;
RAM[16'h06A8] = 8'h00;
RAM[16'h06A9] = 8'h00;
RAM[16'h06AA] = 8'h00;
RAM[16'h06AB] = 8'h00;
RAM[16'h06AC] = 8'h00;
RAM[16'h06AD] = 8'h00;
RAM[16'h06AE] = 8'h00;
RAM[16'h06AF] = 8'h00;
RAM[16'h06B0] = 8'h00;
RAM[16'h06B1] = 8'h00;
RAM[16'h06B2] = 8'h00;
RAM[16'h06B3] = 8'h00;
RAM[16'h06B4] = 8'h00;
RAM[16'h06B5] = 8'h00;
RAM[16'h06B6] = 8'h00;
RAM[16'h06B7] = 8'h00;
RAM[16'h06B8] = 8'h00;
RAM[16'h06B9] = 8'h00;
RAM[16'h06BA] = 8'h00;
RAM[16'h06BB] = 8'h00;
RAM[16'h06BC] = 8'h00;
RAM[16'h06BD] = 8'h00;
RAM[16'h06BE] = 8'h00;
RAM[16'h06BF] = 8'h00;
RAM[16'h06C0] = 8'h00;
RAM[16'h06C1] = 8'h00;
RAM[16'h06C2] = 8'h00;
RAM[16'h06C3] = 8'h00;
RAM[16'h06C4] = 8'h00;
RAM[16'h06C5] = 8'h00;
RAM[16'h06C6] = 8'h00;
RAM[16'h06C7] = 8'h00;
RAM[16'h06C8] = 8'h00;
RAM[16'h06C9] = 8'h00;
RAM[16'h06CA] = 8'h00;
RAM[16'h06CB] = 8'h00;
RAM[16'h06CC] = 8'h00;
RAM[16'h06CD] = 8'h00;
RAM[16'h06CE] = 8'h00;
RAM[16'h06CF] = 8'h00;
RAM[16'h06D0] = 8'h00;
RAM[16'h06D1] = 8'h00;
RAM[16'h06D2] = 8'h00;
RAM[16'h06D3] = 8'h00;
RAM[16'h06D4] = 8'h00;
RAM[16'h06D5] = 8'h00;
RAM[16'h06D6] = 8'h00;
RAM[16'h06D7] = 8'h00;
RAM[16'h06D8] = 8'h00;
RAM[16'h06D9] = 8'h00;
RAM[16'h06DA] = 8'h00;
RAM[16'h06DB] = 8'h00;
RAM[16'h06DC] = 8'h00;
RAM[16'h06DD] = 8'h00;
RAM[16'h06DE] = 8'h00;
RAM[16'h06DF] = 8'h00;
RAM[16'h06E0] = 8'h00;
RAM[16'h06E1] = 8'h00;
RAM[16'h06E2] = 8'h00;
RAM[16'h06E3] = 8'h00;
RAM[16'h06E4] = 8'h00;
RAM[16'h06E5] = 8'h00;
RAM[16'h06E6] = 8'h00;
RAM[16'h06E7] = 8'h00;
RAM[16'h06E8] = 8'h00;
RAM[16'h06E9] = 8'h00;
RAM[16'h06EA] = 8'h00;
RAM[16'h06EB] = 8'h00;
RAM[16'h06EC] = 8'h00;
RAM[16'h06ED] = 8'h00;
RAM[16'h06EE] = 8'h00;
RAM[16'h06EF] = 8'h00;
RAM[16'h06F0] = 8'h00;
RAM[16'h06F1] = 8'h00;
RAM[16'h06F2] = 8'h00;
RAM[16'h06F3] = 8'h00;
RAM[16'h06F4] = 8'h00;
RAM[16'h06F5] = 8'h00;
RAM[16'h06F6] = 8'h00;
RAM[16'h06F7] = 8'h00;
RAM[16'h06F8] = 8'h00;
RAM[16'h06F9] = 8'h00;
RAM[16'h06FA] = 8'h00;
RAM[16'h06FB] = 8'h00;
RAM[16'h06FC] = 8'h00;
RAM[16'h06FD] = 8'h00;
RAM[16'h06FE] = 8'h00;
RAM[16'h06FF] = 8'h00;
RAM[16'h0700] = 8'h00;
RAM[16'h0701] = 8'h00;
RAM[16'h0702] = 8'h00;
RAM[16'h0703] = 8'h00;
RAM[16'h0704] = 8'h00;
RAM[16'h0705] = 8'h00;
RAM[16'h0706] = 8'h00;
RAM[16'h0707] = 8'h00;
RAM[16'h0708] = 8'h00;
RAM[16'h0709] = 8'h00;
RAM[16'h070A] = 8'h00;
RAM[16'h070B] = 8'h00;
RAM[16'h070C] = 8'h00;
RAM[16'h070D] = 8'h00;
RAM[16'h070E] = 8'h00;
RAM[16'h070F] = 8'h00;
RAM[16'h0710] = 8'h00;
RAM[16'h0711] = 8'h00;
RAM[16'h0712] = 8'h00;
RAM[16'h0713] = 8'h00;
RAM[16'h0714] = 8'h00;
RAM[16'h0715] = 8'h00;
RAM[16'h0716] = 8'h00;
RAM[16'h0717] = 8'h00;
RAM[16'h0718] = 8'h00;
RAM[16'h0719] = 8'h00;
RAM[16'h071A] = 8'h00;
RAM[16'h071B] = 8'h00;
RAM[16'h071C] = 8'h00;
RAM[16'h071D] = 8'h00;
RAM[16'h071E] = 8'h00;
RAM[16'h071F] = 8'h00;
RAM[16'h0720] = 8'h00;
RAM[16'h0721] = 8'h00;
RAM[16'h0722] = 8'h00;
RAM[16'h0723] = 8'h00;
RAM[16'h0724] = 8'h00;
RAM[16'h0725] = 8'h00;
RAM[16'h0726] = 8'h00;
RAM[16'h0727] = 8'h00;
RAM[16'h0728] = 8'h00;
RAM[16'h0729] = 8'h00;
RAM[16'h072A] = 8'h00;
RAM[16'h072B] = 8'h00;
RAM[16'h072C] = 8'h00;
RAM[16'h072D] = 8'h00;
RAM[16'h072E] = 8'h00;
RAM[16'h072F] = 8'h00;
RAM[16'h0730] = 8'h00;
RAM[16'h0731] = 8'h00;
RAM[16'h0732] = 8'h00;
RAM[16'h0733] = 8'h00;
RAM[16'h0734] = 8'h00;
RAM[16'h0735] = 8'h00;
RAM[16'h0736] = 8'h00;
RAM[16'h0737] = 8'h00;
RAM[16'h0738] = 8'h00;
RAM[16'h0739] = 8'h00;
RAM[16'h073A] = 8'h00;
RAM[16'h073B] = 8'h00;
RAM[16'h073C] = 8'h00;
RAM[16'h073D] = 8'h00;
RAM[16'h073E] = 8'h00;
RAM[16'h073F] = 8'h00;
RAM[16'h0740] = 8'h00;
RAM[16'h0741] = 8'h00;
RAM[16'h0742] = 8'h00;
RAM[16'h0743] = 8'h00;
RAM[16'h0744] = 8'h00;
RAM[16'h0745] = 8'h00;
RAM[16'h0746] = 8'h00;
RAM[16'h0747] = 8'h00;
RAM[16'h0748] = 8'h00;
RAM[16'h0749] = 8'h00;
RAM[16'h074A] = 8'h00;
RAM[16'h074B] = 8'h00;
RAM[16'h074C] = 8'h00;
RAM[16'h074D] = 8'h00;
RAM[16'h074E] = 8'h00;
RAM[16'h074F] = 8'h00;
RAM[16'h0750] = 8'h00;
RAM[16'h0751] = 8'h00;
RAM[16'h0752] = 8'h00;
RAM[16'h0753] = 8'h00;
RAM[16'h0754] = 8'h00;
RAM[16'h0755] = 8'h00;
RAM[16'h0756] = 8'h00;
RAM[16'h0757] = 8'h00;
RAM[16'h0758] = 8'h00;
RAM[16'h0759] = 8'h00;
RAM[16'h075A] = 8'h00;
RAM[16'h075B] = 8'h00;
RAM[16'h075C] = 8'h00;
RAM[16'h075D] = 8'h00;
RAM[16'h075E] = 8'h00;
RAM[16'h075F] = 8'h00;
RAM[16'h0760] = 8'h00;
RAM[16'h0761] = 8'h00;
RAM[16'h0762] = 8'h00;
RAM[16'h0763] = 8'h00;
RAM[16'h0764] = 8'h00;
RAM[16'h0765] = 8'h00;
RAM[16'h0766] = 8'h00;
RAM[16'h0767] = 8'h00;
RAM[16'h0768] = 8'h00;
RAM[16'h0769] = 8'h00;
RAM[16'h076A] = 8'h00;
RAM[16'h076B] = 8'h00;
RAM[16'h076C] = 8'h00;
RAM[16'h076D] = 8'h00;
RAM[16'h076E] = 8'h00;
RAM[16'h076F] = 8'h00;
RAM[16'h0770] = 8'h00;
RAM[16'h0771] = 8'h00;
RAM[16'h0772] = 8'h00;
RAM[16'h0773] = 8'h00;
RAM[16'h0774] = 8'h00;
RAM[16'h0775] = 8'h00;
RAM[16'h0776] = 8'h00;
RAM[16'h0777] = 8'h00;
RAM[16'h0778] = 8'h00;
RAM[16'h0779] = 8'h00;
RAM[16'h077A] = 8'h00;
RAM[16'h077B] = 8'h00;
RAM[16'h077C] = 8'h00;
RAM[16'h077D] = 8'h00;
RAM[16'h077E] = 8'h00;
RAM[16'h077F] = 8'h00;
RAM[16'h0780] = 8'h00;
RAM[16'h0781] = 8'h00;
RAM[16'h0782] = 8'h00;
RAM[16'h0783] = 8'h00;
RAM[16'h0784] = 8'h00;
RAM[16'h0785] = 8'h00;
RAM[16'h0786] = 8'h00;
RAM[16'h0787] = 8'h00;
RAM[16'h0788] = 8'h00;
RAM[16'h0789] = 8'h00;
RAM[16'h078A] = 8'h00;
RAM[16'h078B] = 8'h00;
RAM[16'h078C] = 8'h00;
RAM[16'h078D] = 8'h00;
RAM[16'h078E] = 8'h00;
RAM[16'h078F] = 8'h00;
RAM[16'h0790] = 8'h00;
RAM[16'h0791] = 8'h00;
RAM[16'h0792] = 8'h00;
RAM[16'h0793] = 8'h00;
RAM[16'h0794] = 8'h00;
RAM[16'h0795] = 8'h00;
RAM[16'h0796] = 8'h00;
RAM[16'h0797] = 8'h00;
RAM[16'h0798] = 8'h00;
RAM[16'h0799] = 8'h00;
RAM[16'h079A] = 8'h00;
RAM[16'h079B] = 8'h00;
RAM[16'h079C] = 8'h00;
RAM[16'h079D] = 8'h00;
RAM[16'h079E] = 8'h00;
RAM[16'h079F] = 8'h00;
RAM[16'h07A0] = 8'h00;
RAM[16'h07A1] = 8'h00;
RAM[16'h07A2] = 8'h00;
RAM[16'h07A3] = 8'h00;
RAM[16'h07A4] = 8'h00;
RAM[16'h07A5] = 8'h00;
RAM[16'h07A6] = 8'h00;
RAM[16'h07A7] = 8'h00;
RAM[16'h07A8] = 8'h00;
RAM[16'h07A9] = 8'h00;
RAM[16'h07AA] = 8'h00;
RAM[16'h07AB] = 8'h00;
RAM[16'h07AC] = 8'h00;
RAM[16'h07AD] = 8'h00;
RAM[16'h07AE] = 8'h00;
RAM[16'h07AF] = 8'h00;
RAM[16'h07B0] = 8'h00;
RAM[16'h07B1] = 8'h00;
RAM[16'h07B2] = 8'h00;
RAM[16'h07B3] = 8'h00;
RAM[16'h07B4] = 8'h00;
RAM[16'h07B5] = 8'h00;
RAM[16'h07B6] = 8'h00;
RAM[16'h07B7] = 8'h00;
RAM[16'h07B8] = 8'h00;
RAM[16'h07B9] = 8'h00;
RAM[16'h07BA] = 8'h00;
RAM[16'h07BB] = 8'h00;
RAM[16'h07BC] = 8'h00;
RAM[16'h07BD] = 8'h00;
RAM[16'h07BE] = 8'h00;
RAM[16'h07BF] = 8'h00;
RAM[16'h07C0] = 8'h00;
RAM[16'h07C1] = 8'h00;
RAM[16'h07C2] = 8'h00;
RAM[16'h07C3] = 8'h00;
RAM[16'h07C4] = 8'h00;
RAM[16'h07C5] = 8'h00;
RAM[16'h07C6] = 8'h00;
RAM[16'h07C7] = 8'h00;
RAM[16'h07C8] = 8'h00;
RAM[16'h07C9] = 8'h00;
RAM[16'h07CA] = 8'h00;
RAM[16'h07CB] = 8'h00;
RAM[16'h07CC] = 8'h00;
RAM[16'h07CD] = 8'h00;
RAM[16'h07CE] = 8'h00;
RAM[16'h07CF] = 8'h00;
RAM[16'h07D0] = 8'h00;
RAM[16'h07D1] = 8'h00;
RAM[16'h07D2] = 8'h00;
RAM[16'h07D3] = 8'h00;
RAM[16'h07D4] = 8'h00;
RAM[16'h07D5] = 8'h00;
RAM[16'h07D6] = 8'h00;
RAM[16'h07D7] = 8'h00;
RAM[16'h07D8] = 8'h00;
RAM[16'h07D9] = 8'h00;
RAM[16'h07DA] = 8'h00;
RAM[16'h07DB] = 8'h00;
RAM[16'h07DC] = 8'h00;
RAM[16'h07DD] = 8'h00;
RAM[16'h07DE] = 8'h00;
RAM[16'h07DF] = 8'h00;
RAM[16'h07E0] = 8'h00;
RAM[16'h07E1] = 8'h00;
RAM[16'h07E2] = 8'h00;
RAM[16'h07E3] = 8'h00;
RAM[16'h07E4] = 8'h00;
RAM[16'h07E5] = 8'h00;
RAM[16'h07E6] = 8'h00;
RAM[16'h07E7] = 8'h00;
RAM[16'h07E8] = 8'h00;
RAM[16'h07E9] = 8'h00;
RAM[16'h07EA] = 8'h00;
RAM[16'h07EB] = 8'h00;
RAM[16'h07EC] = 8'h00;
RAM[16'h07ED] = 8'h00;
RAM[16'h07EE] = 8'h00;
RAM[16'h07EF] = 8'h00;
RAM[16'h07F0] = 8'h00;
RAM[16'h07F1] = 8'h00;
RAM[16'h07F2] = 8'h00;
RAM[16'h07F3] = 8'h00;
RAM[16'h07F4] = 8'h00;
RAM[16'h07F5] = 8'h00;
RAM[16'h07F6] = 8'h00;
RAM[16'h07F7] = 8'h00;
RAM[16'h07F8] = 8'h00;
RAM[16'h07F9] = 8'h00;
RAM[16'h07FA] = 8'h00;
RAM[16'h07FB] = 8'h00;
RAM[16'h07FC] = 8'h00;
RAM[16'h07FD] = 8'h00;
RAM[16'h07FE] = 8'h00;
RAM[16'h07FF] = 8'h00;
RAM[16'h0800] = 8'h00;
RAM[16'h0801] = 8'h00;
RAM[16'h0802] = 8'h00;
RAM[16'h0803] = 8'h00;
RAM[16'h0804] = 8'h00;
RAM[16'h0805] = 8'h00;
RAM[16'h0806] = 8'h00;
RAM[16'h0807] = 8'h00;
RAM[16'h0808] = 8'h00;
RAM[16'h0809] = 8'h00;
RAM[16'h080A] = 8'h00;
RAM[16'h080B] = 8'h00;
RAM[16'h080C] = 8'h00;
RAM[16'h080D] = 8'h00;
RAM[16'h080E] = 8'h00;
RAM[16'h080F] = 8'h00;
RAM[16'h0810] = 8'h00;
RAM[16'h0811] = 8'h00;
RAM[16'h0812] = 8'h00;
RAM[16'h0813] = 8'h00;
RAM[16'h0814] = 8'h00;
RAM[16'h0815] = 8'h00;
RAM[16'h0816] = 8'h00;
RAM[16'h0817] = 8'h00;
RAM[16'h0818] = 8'h00;
RAM[16'h0819] = 8'h00;
RAM[16'h081A] = 8'h00;
RAM[16'h081B] = 8'h00;
RAM[16'h081C] = 8'h00;
RAM[16'h081D] = 8'h00;
RAM[16'h081E] = 8'h00;
RAM[16'h081F] = 8'h00;
RAM[16'h0820] = 8'h00;
RAM[16'h0821] = 8'h00;
RAM[16'h0822] = 8'h00;
RAM[16'h0823] = 8'h00;
RAM[16'h0824] = 8'h00;
RAM[16'h0825] = 8'h00;
RAM[16'h0826] = 8'h00;
RAM[16'h0827] = 8'h00;
RAM[16'h0828] = 8'h00;
RAM[16'h0829] = 8'h00;
RAM[16'h082A] = 8'h00;
RAM[16'h082B] = 8'h00;
RAM[16'h082C] = 8'h00;
RAM[16'h082D] = 8'h00;
RAM[16'h082E] = 8'h00;
RAM[16'h082F] = 8'h00;
RAM[16'h0830] = 8'h00;
RAM[16'h0831] = 8'h00;
RAM[16'h0832] = 8'h00;
RAM[16'h0833] = 8'h00;
RAM[16'h0834] = 8'h00;
RAM[16'h0835] = 8'h00;
RAM[16'h0836] = 8'h00;
RAM[16'h0837] = 8'h00;
RAM[16'h0838] = 8'h00;
RAM[16'h0839] = 8'h00;
RAM[16'h083A] = 8'h00;
RAM[16'h083B] = 8'h00;
RAM[16'h083C] = 8'h00;
RAM[16'h083D] = 8'h00;
RAM[16'h083E] = 8'h00;
RAM[16'h083F] = 8'h00;
RAM[16'h0840] = 8'h00;
RAM[16'h0841] = 8'h00;
RAM[16'h0842] = 8'h00;
RAM[16'h0843] = 8'h00;
RAM[16'h0844] = 8'h00;
RAM[16'h0845] = 8'h00;
RAM[16'h0846] = 8'h00;
RAM[16'h0847] = 8'h00;
RAM[16'h0848] = 8'h00;
RAM[16'h0849] = 8'h00;
RAM[16'h084A] = 8'h00;
RAM[16'h084B] = 8'h00;
RAM[16'h084C] = 8'h00;
RAM[16'h084D] = 8'h00;
RAM[16'h084E] = 8'h00;
RAM[16'h084F] = 8'h00;
RAM[16'h0850] = 8'h00;
RAM[16'h0851] = 8'h00;
RAM[16'h0852] = 8'h00;
RAM[16'h0853] = 8'h00;
RAM[16'h0854] = 8'h00;
RAM[16'h0855] = 8'h00;
RAM[16'h0856] = 8'h00;
RAM[16'h0857] = 8'h00;
RAM[16'h0858] = 8'h00;
RAM[16'h0859] = 8'h00;
RAM[16'h085A] = 8'h00;
RAM[16'h085B] = 8'h00;
RAM[16'h085C] = 8'h00;
RAM[16'h085D] = 8'h00;
RAM[16'h085E] = 8'h00;
RAM[16'h085F] = 8'h00;
RAM[16'h0860] = 8'h00;
RAM[16'h0861] = 8'h00;
RAM[16'h0862] = 8'h00;
RAM[16'h0863] = 8'h00;
RAM[16'h0864] = 8'h00;
RAM[16'h0865] = 8'h00;
RAM[16'h0866] = 8'h00;
RAM[16'h0867] = 8'h00;
RAM[16'h0868] = 8'h00;
RAM[16'h0869] = 8'h00;
RAM[16'h086A] = 8'h00;
RAM[16'h086B] = 8'h00;
RAM[16'h086C] = 8'h00;
RAM[16'h086D] = 8'h00;
RAM[16'h086E] = 8'h00;
RAM[16'h086F] = 8'h00;
RAM[16'h0870] = 8'h00;
RAM[16'h0871] = 8'h00;
RAM[16'h0872] = 8'h00;
RAM[16'h0873] = 8'h00;
RAM[16'h0874] = 8'h00;
RAM[16'h0875] = 8'h00;
RAM[16'h0876] = 8'h00;
RAM[16'h0877] = 8'h00;
RAM[16'h0878] = 8'h00;
RAM[16'h0879] = 8'h00;
RAM[16'h087A] = 8'h00;
RAM[16'h087B] = 8'h00;
RAM[16'h087C] = 8'h00;
RAM[16'h087D] = 8'h00;
RAM[16'h087E] = 8'h00;
RAM[16'h087F] = 8'h00;
RAM[16'h0880] = 8'h00;
RAM[16'h0881] = 8'h00;
RAM[16'h0882] = 8'h00;
RAM[16'h0883] = 8'h00;
RAM[16'h0884] = 8'h00;
RAM[16'h0885] = 8'h00;
RAM[16'h0886] = 8'h00;
RAM[16'h0887] = 8'h00;
RAM[16'h0888] = 8'h00;
RAM[16'h0889] = 8'h00;
RAM[16'h088A] = 8'h00;
RAM[16'h088B] = 8'h00;
RAM[16'h088C] = 8'h00;
RAM[16'h088D] = 8'h00;
RAM[16'h088E] = 8'h00;
RAM[16'h088F] = 8'h00;
RAM[16'h0890] = 8'h00;
RAM[16'h0891] = 8'h00;
RAM[16'h0892] = 8'h00;
RAM[16'h0893] = 8'h00;
RAM[16'h0894] = 8'h00;
RAM[16'h0895] = 8'h00;
RAM[16'h0896] = 8'h00;
RAM[16'h0897] = 8'h00;
RAM[16'h0898] = 8'h00;
RAM[16'h0899] = 8'h00;
RAM[16'h089A] = 8'h00;
RAM[16'h089B] = 8'h00;
RAM[16'h089C] = 8'h00;
RAM[16'h089D] = 8'h00;
RAM[16'h089E] = 8'h00;
RAM[16'h089F] = 8'h00;
RAM[16'h08A0] = 8'h00;
RAM[16'h08A1] = 8'h00;
RAM[16'h08A2] = 8'h00;
RAM[16'h08A3] = 8'h00;
RAM[16'h08A4] = 8'h00;
RAM[16'h08A5] = 8'h00;
RAM[16'h08A6] = 8'h00;
RAM[16'h08A7] = 8'h00;
RAM[16'h08A8] = 8'h00;
RAM[16'h08A9] = 8'h00;
RAM[16'h08AA] = 8'h00;
RAM[16'h08AB] = 8'h00;
RAM[16'h08AC] = 8'h00;
RAM[16'h08AD] = 8'h00;
RAM[16'h08AE] = 8'h00;
RAM[16'h08AF] = 8'h00;
RAM[16'h08B0] = 8'h00;
RAM[16'h08B1] = 8'h00;
RAM[16'h08B2] = 8'h00;
RAM[16'h08B3] = 8'h00;
RAM[16'h08B4] = 8'h00;
RAM[16'h08B5] = 8'h00;
RAM[16'h08B6] = 8'h00;
RAM[16'h08B7] = 8'h00;
RAM[16'h08B8] = 8'h00;
RAM[16'h08B9] = 8'h00;
RAM[16'h08BA] = 8'h00;
RAM[16'h08BB] = 8'h00;
RAM[16'h08BC] = 8'h00;
RAM[16'h08BD] = 8'h00;
RAM[16'h08BE] = 8'h00;
RAM[16'h08BF] = 8'h00;
RAM[16'h08C0] = 8'h00;
RAM[16'h08C1] = 8'h00;
RAM[16'h08C2] = 8'h00;
RAM[16'h08C3] = 8'h00;
RAM[16'h08C4] = 8'h00;
RAM[16'h08C5] = 8'h00;
RAM[16'h08C6] = 8'h00;
RAM[16'h08C7] = 8'h00;
RAM[16'h08C8] = 8'h00;
RAM[16'h08C9] = 8'h00;
RAM[16'h08CA] = 8'h00;
RAM[16'h08CB] = 8'h00;
RAM[16'h08CC] = 8'h00;
RAM[16'h08CD] = 8'h00;
RAM[16'h08CE] = 8'h00;
RAM[16'h08CF] = 8'h00;
RAM[16'h08D0] = 8'h00;
RAM[16'h08D1] = 8'h00;
RAM[16'h08D2] = 8'h00;
RAM[16'h08D3] = 8'h00;
RAM[16'h08D4] = 8'h00;
RAM[16'h08D5] = 8'h00;
RAM[16'h08D6] = 8'h00;
RAM[16'h08D7] = 8'h00;
RAM[16'h08D8] = 8'h00;
RAM[16'h08D9] = 8'h00;
RAM[16'h08DA] = 8'h00;
RAM[16'h08DB] = 8'h00;
RAM[16'h08DC] = 8'h00;
RAM[16'h08DD] = 8'h00;
RAM[16'h08DE] = 8'h00;
RAM[16'h08DF] = 8'h00;
RAM[16'h08E0] = 8'h00;
RAM[16'h08E1] = 8'h00;
RAM[16'h08E2] = 8'h00;
RAM[16'h08E3] = 8'h00;
RAM[16'h08E4] = 8'h00;
RAM[16'h08E5] = 8'h00;
RAM[16'h08E6] = 8'h00;
RAM[16'h08E7] = 8'h00;
RAM[16'h08E8] = 8'h00;
RAM[16'h08E9] = 8'h00;
RAM[16'h08EA] = 8'h00;
RAM[16'h08EB] = 8'h00;
RAM[16'h08EC] = 8'h00;
RAM[16'h08ED] = 8'h00;
RAM[16'h08EE] = 8'h00;
RAM[16'h08EF] = 8'h00;
RAM[16'h08F0] = 8'h00;
RAM[16'h08F1] = 8'h00;
RAM[16'h08F2] = 8'h00;
RAM[16'h08F3] = 8'h00;
RAM[16'h08F4] = 8'h00;
RAM[16'h08F5] = 8'h00;
RAM[16'h08F6] = 8'h00;
RAM[16'h08F7] = 8'h00;
RAM[16'h08F8] = 8'h00;
RAM[16'h08F9] = 8'h00;
RAM[16'h08FA] = 8'h00;
RAM[16'h08FB] = 8'h00;
RAM[16'h08FC] = 8'h00;
RAM[16'h08FD] = 8'h00;
RAM[16'h08FE] = 8'h00;
RAM[16'h08FF] = 8'h00;
RAM[16'h0900] = 8'h00;
RAM[16'h0901] = 8'h00;
RAM[16'h0902] = 8'h00;
RAM[16'h0903] = 8'h00;
RAM[16'h0904] = 8'h00;
RAM[16'h0905] = 8'h00;
RAM[16'h0906] = 8'h00;
RAM[16'h0907] = 8'h00;
RAM[16'h0908] = 8'h00;
RAM[16'h0909] = 8'h00;
RAM[16'h090A] = 8'h00;
RAM[16'h090B] = 8'h00;
RAM[16'h090C] = 8'h00;
RAM[16'h090D] = 8'h00;
RAM[16'h090E] = 8'h00;
RAM[16'h090F] = 8'h00;
RAM[16'h0910] = 8'h00;
RAM[16'h0911] = 8'h00;
RAM[16'h0912] = 8'h00;
RAM[16'h0913] = 8'h00;
RAM[16'h0914] = 8'h00;
RAM[16'h0915] = 8'h00;
RAM[16'h0916] = 8'h00;
RAM[16'h0917] = 8'h00;
RAM[16'h0918] = 8'h00;
RAM[16'h0919] = 8'h00;
RAM[16'h091A] = 8'h00;
RAM[16'h091B] = 8'h00;
RAM[16'h091C] = 8'h00;
RAM[16'h091D] = 8'h00;
RAM[16'h091E] = 8'h00;
RAM[16'h091F] = 8'h00;
RAM[16'h0920] = 8'h00;
RAM[16'h0921] = 8'h00;
RAM[16'h0922] = 8'h00;
RAM[16'h0923] = 8'h00;
RAM[16'h0924] = 8'h00;
RAM[16'h0925] = 8'h00;
RAM[16'h0926] = 8'h00;
RAM[16'h0927] = 8'h00;
RAM[16'h0928] = 8'h00;
RAM[16'h0929] = 8'h00;
RAM[16'h092A] = 8'h00;
RAM[16'h092B] = 8'h00;
RAM[16'h092C] = 8'h00;
RAM[16'h092D] = 8'h00;
RAM[16'h092E] = 8'h00;
RAM[16'h092F] = 8'h00;
RAM[16'h0930] = 8'h00;
RAM[16'h0931] = 8'h00;
RAM[16'h0932] = 8'h00;
RAM[16'h0933] = 8'h00;
RAM[16'h0934] = 8'h00;
RAM[16'h0935] = 8'h00;
RAM[16'h0936] = 8'h00;
RAM[16'h0937] = 8'h00;
RAM[16'h0938] = 8'h00;
RAM[16'h0939] = 8'h00;
RAM[16'h093A] = 8'h00;
RAM[16'h093B] = 8'h00;
RAM[16'h093C] = 8'h00;
RAM[16'h093D] = 8'h00;
RAM[16'h093E] = 8'h00;
RAM[16'h093F] = 8'h00;
RAM[16'h0940] = 8'h00;
RAM[16'h0941] = 8'h00;
RAM[16'h0942] = 8'h00;
RAM[16'h0943] = 8'h00;
RAM[16'h0944] = 8'h00;
RAM[16'h0945] = 8'h00;
RAM[16'h0946] = 8'h00;
RAM[16'h0947] = 8'h00;
RAM[16'h0948] = 8'h00;
RAM[16'h0949] = 8'h00;
RAM[16'h094A] = 8'h00;
RAM[16'h094B] = 8'h00;
RAM[16'h094C] = 8'h00;
RAM[16'h094D] = 8'h00;
RAM[16'h094E] = 8'h00;
RAM[16'h094F] = 8'h00;
RAM[16'h0950] = 8'h00;
RAM[16'h0951] = 8'h00;
RAM[16'h0952] = 8'h00;
RAM[16'h0953] = 8'h00;
RAM[16'h0954] = 8'h00;
RAM[16'h0955] = 8'h00;
RAM[16'h0956] = 8'h00;
RAM[16'h0957] = 8'h00;
RAM[16'h0958] = 8'h00;
RAM[16'h0959] = 8'h00;
RAM[16'h095A] = 8'h00;
RAM[16'h095B] = 8'h00;
RAM[16'h095C] = 8'h00;
RAM[16'h095D] = 8'h00;
RAM[16'h095E] = 8'h00;
RAM[16'h095F] = 8'h00;
RAM[16'h0960] = 8'h00;
RAM[16'h0961] = 8'h00;
RAM[16'h0962] = 8'h00;
RAM[16'h0963] = 8'h00;
RAM[16'h0964] = 8'h00;
RAM[16'h0965] = 8'h00;
RAM[16'h0966] = 8'h00;
RAM[16'h0967] = 8'h00;
RAM[16'h0968] = 8'h00;
RAM[16'h0969] = 8'h00;
RAM[16'h096A] = 8'h00;
RAM[16'h096B] = 8'h00;
RAM[16'h096C] = 8'h00;
RAM[16'h096D] = 8'h00;
RAM[16'h096E] = 8'h00;
RAM[16'h096F] = 8'h00;
RAM[16'h0970] = 8'h00;
RAM[16'h0971] = 8'h00;
RAM[16'h0972] = 8'h00;
RAM[16'h0973] = 8'h00;
RAM[16'h0974] = 8'h00;
RAM[16'h0975] = 8'h00;
RAM[16'h0976] = 8'h00;
RAM[16'h0977] = 8'h00;
RAM[16'h0978] = 8'h00;
RAM[16'h0979] = 8'h00;
RAM[16'h097A] = 8'h00;
RAM[16'h097B] = 8'h00;
RAM[16'h097C] = 8'h00;
RAM[16'h097D] = 8'h00;
RAM[16'h097E] = 8'h00;
RAM[16'h097F] = 8'h00;
RAM[16'h0980] = 8'h00;
RAM[16'h0981] = 8'h00;
RAM[16'h0982] = 8'h00;
RAM[16'h0983] = 8'h00;
RAM[16'h0984] = 8'h00;
RAM[16'h0985] = 8'h00;
RAM[16'h0986] = 8'h00;
RAM[16'h0987] = 8'h00;
RAM[16'h0988] = 8'h00;
RAM[16'h0989] = 8'h00;
RAM[16'h098A] = 8'h00;
RAM[16'h098B] = 8'h00;
RAM[16'h098C] = 8'h00;
RAM[16'h098D] = 8'h00;
RAM[16'h098E] = 8'h00;
RAM[16'h098F] = 8'h00;
RAM[16'h0990] = 8'h00;
RAM[16'h0991] = 8'h00;
RAM[16'h0992] = 8'h00;
RAM[16'h0993] = 8'h00;
RAM[16'h0994] = 8'h00;
RAM[16'h0995] = 8'h00;
RAM[16'h0996] = 8'h00;
RAM[16'h0997] = 8'h00;
RAM[16'h0998] = 8'h00;
RAM[16'h0999] = 8'h00;
RAM[16'h099A] = 8'h00;
RAM[16'h099B] = 8'h00;
RAM[16'h099C] = 8'h00;
RAM[16'h099D] = 8'h00;
RAM[16'h099E] = 8'h00;
RAM[16'h099F] = 8'h00;
RAM[16'h09A0] = 8'h00;
RAM[16'h09A1] = 8'h00;
RAM[16'h09A2] = 8'h00;
RAM[16'h09A3] = 8'h00;
RAM[16'h09A4] = 8'h00;
RAM[16'h09A5] = 8'h00;
RAM[16'h09A6] = 8'h00;
RAM[16'h09A7] = 8'h00;
RAM[16'h09A8] = 8'h00;
RAM[16'h09A9] = 8'h00;
RAM[16'h09AA] = 8'h00;
RAM[16'h09AB] = 8'h00;
RAM[16'h09AC] = 8'h00;
RAM[16'h09AD] = 8'h00;
RAM[16'h09AE] = 8'h00;
RAM[16'h09AF] = 8'h00;
RAM[16'h09B0] = 8'h00;
RAM[16'h09B1] = 8'h00;
RAM[16'h09B2] = 8'h00;
RAM[16'h09B3] = 8'h00;
RAM[16'h09B4] = 8'h00;
RAM[16'h09B5] = 8'h00;
RAM[16'h09B6] = 8'h00;
RAM[16'h09B7] = 8'h00;
RAM[16'h09B8] = 8'h00;
RAM[16'h09B9] = 8'h00;
RAM[16'h09BA] = 8'h00;
RAM[16'h09BB] = 8'h00;
RAM[16'h09BC] = 8'h00;
RAM[16'h09BD] = 8'h00;
RAM[16'h09BE] = 8'h00;
RAM[16'h09BF] = 8'h00;
RAM[16'h09C0] = 8'h00;
RAM[16'h09C1] = 8'h00;
RAM[16'h09C2] = 8'h00;
RAM[16'h09C3] = 8'h00;
RAM[16'h09C4] = 8'h00;
RAM[16'h09C5] = 8'h00;
RAM[16'h09C6] = 8'h00;
RAM[16'h09C7] = 8'h00;
RAM[16'h09C8] = 8'h00;
RAM[16'h09C9] = 8'h00;
RAM[16'h09CA] = 8'h00;
RAM[16'h09CB] = 8'h00;
RAM[16'h09CC] = 8'h00;
RAM[16'h09CD] = 8'h00;
RAM[16'h09CE] = 8'h00;
RAM[16'h09CF] = 8'h00;
RAM[16'h09D0] = 8'h00;
RAM[16'h09D1] = 8'h00;
RAM[16'h09D2] = 8'h00;
RAM[16'h09D3] = 8'h00;
RAM[16'h09D4] = 8'h00;
RAM[16'h09D5] = 8'h00;
RAM[16'h09D6] = 8'h00;
RAM[16'h09D7] = 8'h00;
RAM[16'h09D8] = 8'h00;
RAM[16'h09D9] = 8'h00;
RAM[16'h09DA] = 8'h00;
RAM[16'h09DB] = 8'h00;
RAM[16'h09DC] = 8'h00;
RAM[16'h09DD] = 8'h00;
RAM[16'h09DE] = 8'h00;
RAM[16'h09DF] = 8'h00;
RAM[16'h09E0] = 8'h00;
RAM[16'h09E1] = 8'h00;
RAM[16'h09E2] = 8'h00;
RAM[16'h09E3] = 8'h00;
RAM[16'h09E4] = 8'h00;
RAM[16'h09E5] = 8'h00;
RAM[16'h09E6] = 8'h00;
RAM[16'h09E7] = 8'h00;
RAM[16'h09E8] = 8'h00;
RAM[16'h09E9] = 8'h00;
RAM[16'h09EA] = 8'h00;
RAM[16'h09EB] = 8'h00;
RAM[16'h09EC] = 8'h00;
RAM[16'h09ED] = 8'h00;
RAM[16'h09EE] = 8'h00;
RAM[16'h09EF] = 8'h00;
RAM[16'h09F0] = 8'h00;
RAM[16'h09F1] = 8'h00;
RAM[16'h09F2] = 8'h00;
RAM[16'h09F3] = 8'h00;
RAM[16'h09F4] = 8'h00;
RAM[16'h09F5] = 8'h00;
RAM[16'h09F6] = 8'h00;
RAM[16'h09F7] = 8'h00;
RAM[16'h09F8] = 8'h00;
RAM[16'h09F9] = 8'h00;
RAM[16'h09FA] = 8'h00;
RAM[16'h09FB] = 8'h00;
RAM[16'h09FC] = 8'h00;
RAM[16'h09FD] = 8'h00;
RAM[16'h09FE] = 8'h00;
RAM[16'h09FF] = 8'h00;
RAM[16'h0A00] = 8'h00;
RAM[16'h0A01] = 8'h00;
RAM[16'h0A02] = 8'h00;
RAM[16'h0A03] = 8'h00;
RAM[16'h0A04] = 8'h00;
RAM[16'h0A05] = 8'h00;
RAM[16'h0A06] = 8'h00;
RAM[16'h0A07] = 8'h00;
RAM[16'h0A08] = 8'h00;
RAM[16'h0A09] = 8'h00;
RAM[16'h0A0A] = 8'h00;
RAM[16'h0A0B] = 8'h00;
RAM[16'h0A0C] = 8'h00;
RAM[16'h0A0D] = 8'h00;
RAM[16'h0A0E] = 8'h00;
RAM[16'h0A0F] = 8'h00;
RAM[16'h0A10] = 8'h00;
RAM[16'h0A11] = 8'h00;
RAM[16'h0A12] = 8'h00;
RAM[16'h0A13] = 8'h00;
RAM[16'h0A14] = 8'h00;
RAM[16'h0A15] = 8'h00;
RAM[16'h0A16] = 8'h00;
RAM[16'h0A17] = 8'h00;
RAM[16'h0A18] = 8'h00;
RAM[16'h0A19] = 8'h00;
RAM[16'h0A1A] = 8'h00;
RAM[16'h0A1B] = 8'h00;
RAM[16'h0A1C] = 8'h00;
RAM[16'h0A1D] = 8'h00;
RAM[16'h0A1E] = 8'h00;
RAM[16'h0A1F] = 8'h00;
RAM[16'h0A20] = 8'h00;
RAM[16'h0A21] = 8'h00;
RAM[16'h0A22] = 8'h00;
RAM[16'h0A23] = 8'h00;
RAM[16'h0A24] = 8'h00;
RAM[16'h0A25] = 8'h00;
RAM[16'h0A26] = 8'h00;
RAM[16'h0A27] = 8'h00;
RAM[16'h0A28] = 8'h00;
RAM[16'h0A29] = 8'h00;
RAM[16'h0A2A] = 8'h00;
RAM[16'h0A2B] = 8'h00;
RAM[16'h0A2C] = 8'h00;
RAM[16'h0A2D] = 8'h00;
RAM[16'h0A2E] = 8'h00;
RAM[16'h0A2F] = 8'h00;
RAM[16'h0A30] = 8'h00;
RAM[16'h0A31] = 8'h00;
RAM[16'h0A32] = 8'h00;
RAM[16'h0A33] = 8'h00;
RAM[16'h0A34] = 8'h00;
RAM[16'h0A35] = 8'h00;
RAM[16'h0A36] = 8'h00;
RAM[16'h0A37] = 8'h00;
RAM[16'h0A38] = 8'h00;
RAM[16'h0A39] = 8'h00;
RAM[16'h0A3A] = 8'h00;
RAM[16'h0A3B] = 8'h00;
RAM[16'h0A3C] = 8'h00;
RAM[16'h0A3D] = 8'h00;
RAM[16'h0A3E] = 8'h00;
RAM[16'h0A3F] = 8'h00;
RAM[16'h0A40] = 8'h00;
RAM[16'h0A41] = 8'h00;
RAM[16'h0A42] = 8'h00;
RAM[16'h0A43] = 8'h00;
RAM[16'h0A44] = 8'h00;
RAM[16'h0A45] = 8'h00;
RAM[16'h0A46] = 8'h00;
RAM[16'h0A47] = 8'h00;
RAM[16'h0A48] = 8'h00;
RAM[16'h0A49] = 8'h00;
RAM[16'h0A4A] = 8'h00;
RAM[16'h0A4B] = 8'h00;
RAM[16'h0A4C] = 8'h00;
RAM[16'h0A4D] = 8'h00;
RAM[16'h0A4E] = 8'h00;
RAM[16'h0A4F] = 8'h00;
RAM[16'h0A50] = 8'h00;
RAM[16'h0A51] = 8'h00;
RAM[16'h0A52] = 8'h00;
RAM[16'h0A53] = 8'h00;
RAM[16'h0A54] = 8'h00;
RAM[16'h0A55] = 8'h00;
RAM[16'h0A56] = 8'h00;
RAM[16'h0A57] = 8'h00;
RAM[16'h0A58] = 8'h00;
RAM[16'h0A59] = 8'h00;
RAM[16'h0A5A] = 8'h00;
RAM[16'h0A5B] = 8'h00;
RAM[16'h0A5C] = 8'h00;
RAM[16'h0A5D] = 8'h00;
RAM[16'h0A5E] = 8'h00;
RAM[16'h0A5F] = 8'h00;
RAM[16'h0A60] = 8'h00;
RAM[16'h0A61] = 8'h00;
RAM[16'h0A62] = 8'h00;
RAM[16'h0A63] = 8'h00;
RAM[16'h0A64] = 8'h00;
RAM[16'h0A65] = 8'h00;
RAM[16'h0A66] = 8'h00;
RAM[16'h0A67] = 8'h00;
RAM[16'h0A68] = 8'h00;
RAM[16'h0A69] = 8'h00;
RAM[16'h0A6A] = 8'h00;
RAM[16'h0A6B] = 8'h00;
RAM[16'h0A6C] = 8'h00;
RAM[16'h0A6D] = 8'h00;
RAM[16'h0A6E] = 8'h00;
RAM[16'h0A6F] = 8'h00;
RAM[16'h0A70] = 8'h00;
RAM[16'h0A71] = 8'h00;
RAM[16'h0A72] = 8'h00;
RAM[16'h0A73] = 8'h00;
RAM[16'h0A74] = 8'h00;
RAM[16'h0A75] = 8'h00;
RAM[16'h0A76] = 8'h00;
RAM[16'h0A77] = 8'h00;
RAM[16'h0A78] = 8'h00;
RAM[16'h0A79] = 8'h00;
RAM[16'h0A7A] = 8'h00;
RAM[16'h0A7B] = 8'h00;
RAM[16'h0A7C] = 8'h00;
RAM[16'h0A7D] = 8'h00;
RAM[16'h0A7E] = 8'h00;
RAM[16'h0A7F] = 8'h00;
RAM[16'h0A80] = 8'h00;
RAM[16'h0A81] = 8'h00;
RAM[16'h0A82] = 8'h00;
RAM[16'h0A83] = 8'h00;
RAM[16'h0A84] = 8'h00;
RAM[16'h0A85] = 8'h00;
RAM[16'h0A86] = 8'h00;
RAM[16'h0A87] = 8'h00;
RAM[16'h0A88] = 8'h00;
RAM[16'h0A89] = 8'h00;
RAM[16'h0A8A] = 8'h00;
RAM[16'h0A8B] = 8'h00;
RAM[16'h0A8C] = 8'h00;
RAM[16'h0A8D] = 8'h00;
RAM[16'h0A8E] = 8'h00;
RAM[16'h0A8F] = 8'h00;
RAM[16'h0A90] = 8'h00;
RAM[16'h0A91] = 8'h00;
RAM[16'h0A92] = 8'h00;
RAM[16'h0A93] = 8'h00;
RAM[16'h0A94] = 8'h00;
RAM[16'h0A95] = 8'h00;
RAM[16'h0A96] = 8'h00;
RAM[16'h0A97] = 8'h00;
RAM[16'h0A98] = 8'h00;
RAM[16'h0A99] = 8'h00;
RAM[16'h0A9A] = 8'h00;
RAM[16'h0A9B] = 8'h00;
RAM[16'h0A9C] = 8'h00;
RAM[16'h0A9D] = 8'h00;
RAM[16'h0A9E] = 8'h00;
RAM[16'h0A9F] = 8'h00;
RAM[16'h0AA0] = 8'h00;
RAM[16'h0AA1] = 8'h00;
RAM[16'h0AA2] = 8'h00;
RAM[16'h0AA3] = 8'h00;
RAM[16'h0AA4] = 8'h00;
RAM[16'h0AA5] = 8'h00;
RAM[16'h0AA6] = 8'h00;
RAM[16'h0AA7] = 8'h00;
RAM[16'h0AA8] = 8'h00;
RAM[16'h0AA9] = 8'h00;
RAM[16'h0AAA] = 8'h00;
RAM[16'h0AAB] = 8'h00;
RAM[16'h0AAC] = 8'h00;
RAM[16'h0AAD] = 8'h00;
RAM[16'h0AAE] = 8'h00;
RAM[16'h0AAF] = 8'h00;
RAM[16'h0AB0] = 8'h00;
RAM[16'h0AB1] = 8'h00;
RAM[16'h0AB2] = 8'h00;
RAM[16'h0AB3] = 8'h00;
RAM[16'h0AB4] = 8'h00;
RAM[16'h0AB5] = 8'h00;
RAM[16'h0AB6] = 8'h00;
RAM[16'h0AB7] = 8'h00;
RAM[16'h0AB8] = 8'h00;
RAM[16'h0AB9] = 8'h00;
RAM[16'h0ABA] = 8'h00;
RAM[16'h0ABB] = 8'h00;
RAM[16'h0ABC] = 8'h00;
RAM[16'h0ABD] = 8'h00;
RAM[16'h0ABE] = 8'h00;
RAM[16'h0ABF] = 8'h00;
RAM[16'h0AC0] = 8'h00;
RAM[16'h0AC1] = 8'h00;
RAM[16'h0AC2] = 8'h00;
RAM[16'h0AC3] = 8'h00;
RAM[16'h0AC4] = 8'h00;
RAM[16'h0AC5] = 8'h00;
RAM[16'h0AC6] = 8'h00;
RAM[16'h0AC7] = 8'h00;
RAM[16'h0AC8] = 8'h00;
RAM[16'h0AC9] = 8'h00;
RAM[16'h0ACA] = 8'h00;
RAM[16'h0ACB] = 8'h00;
RAM[16'h0ACC] = 8'h00;
RAM[16'h0ACD] = 8'h00;
RAM[16'h0ACE] = 8'h00;
RAM[16'h0ACF] = 8'h00;
RAM[16'h0AD0] = 8'h00;
RAM[16'h0AD1] = 8'h00;
RAM[16'h0AD2] = 8'h00;
RAM[16'h0AD3] = 8'h00;
RAM[16'h0AD4] = 8'h00;
RAM[16'h0AD5] = 8'h00;
RAM[16'h0AD6] = 8'h00;
RAM[16'h0AD7] = 8'h00;
RAM[16'h0AD8] = 8'h00;
RAM[16'h0AD9] = 8'h00;
RAM[16'h0ADA] = 8'h00;
RAM[16'h0ADB] = 8'h00;
RAM[16'h0ADC] = 8'h00;
RAM[16'h0ADD] = 8'h00;
RAM[16'h0ADE] = 8'h00;
RAM[16'h0ADF] = 8'h00;
RAM[16'h0AE0] = 8'h00;
RAM[16'h0AE1] = 8'h00;
RAM[16'h0AE2] = 8'h00;
RAM[16'h0AE3] = 8'h00;
RAM[16'h0AE4] = 8'h00;
RAM[16'h0AE5] = 8'h00;
RAM[16'h0AE6] = 8'h00;
RAM[16'h0AE7] = 8'h00;
RAM[16'h0AE8] = 8'h00;
RAM[16'h0AE9] = 8'h00;
RAM[16'h0AEA] = 8'h00;
RAM[16'h0AEB] = 8'h00;
RAM[16'h0AEC] = 8'h00;
RAM[16'h0AED] = 8'h00;
RAM[16'h0AEE] = 8'h00;
RAM[16'h0AEF] = 8'h00;
RAM[16'h0AF0] = 8'h00;
RAM[16'h0AF1] = 8'h00;
RAM[16'h0AF2] = 8'h00;
RAM[16'h0AF3] = 8'h00;
RAM[16'h0AF4] = 8'h00;
RAM[16'h0AF5] = 8'h00;
RAM[16'h0AF6] = 8'h00;
RAM[16'h0AF7] = 8'h00;
RAM[16'h0AF8] = 8'h00;
RAM[16'h0AF9] = 8'h00;
RAM[16'h0AFA] = 8'h00;
RAM[16'h0AFB] = 8'h00;
RAM[16'h0AFC] = 8'h00;
RAM[16'h0AFD] = 8'h00;
RAM[16'h0AFE] = 8'h00;
RAM[16'h0AFF] = 8'h00;
RAM[16'h0B00] = 8'h00;
RAM[16'h0B01] = 8'h00;
RAM[16'h0B02] = 8'h00;
RAM[16'h0B03] = 8'h00;
RAM[16'h0B04] = 8'h00;
RAM[16'h0B05] = 8'h00;
RAM[16'h0B06] = 8'h00;
RAM[16'h0B07] = 8'h00;
RAM[16'h0B08] = 8'h00;
RAM[16'h0B09] = 8'h00;
RAM[16'h0B0A] = 8'h00;
RAM[16'h0B0B] = 8'h00;
RAM[16'h0B0C] = 8'h00;
RAM[16'h0B0D] = 8'h00;
RAM[16'h0B0E] = 8'h00;
RAM[16'h0B0F] = 8'h00;
RAM[16'h0B10] = 8'h00;
RAM[16'h0B11] = 8'h00;
RAM[16'h0B12] = 8'h00;
RAM[16'h0B13] = 8'h00;
RAM[16'h0B14] = 8'h00;
RAM[16'h0B15] = 8'h00;
RAM[16'h0B16] = 8'h00;
RAM[16'h0B17] = 8'h00;
RAM[16'h0B18] = 8'h00;
RAM[16'h0B19] = 8'h00;
RAM[16'h0B1A] = 8'h00;
RAM[16'h0B1B] = 8'h00;
RAM[16'h0B1C] = 8'h00;
RAM[16'h0B1D] = 8'h00;
RAM[16'h0B1E] = 8'h00;
RAM[16'h0B1F] = 8'h00;
RAM[16'h0B20] = 8'h00;
RAM[16'h0B21] = 8'h00;
RAM[16'h0B22] = 8'h00;
RAM[16'h0B23] = 8'h00;
RAM[16'h0B24] = 8'h00;
RAM[16'h0B25] = 8'h00;
RAM[16'h0B26] = 8'h00;
RAM[16'h0B27] = 8'h00;
RAM[16'h0B28] = 8'h00;
RAM[16'h0B29] = 8'h00;
RAM[16'h0B2A] = 8'h00;
RAM[16'h0B2B] = 8'h00;
RAM[16'h0B2C] = 8'h00;
RAM[16'h0B2D] = 8'h00;
RAM[16'h0B2E] = 8'h00;
RAM[16'h0B2F] = 8'h00;
RAM[16'h0B30] = 8'h00;
RAM[16'h0B31] = 8'h00;
RAM[16'h0B32] = 8'h00;
RAM[16'h0B33] = 8'h00;
RAM[16'h0B34] = 8'h00;
RAM[16'h0B35] = 8'h00;
RAM[16'h0B36] = 8'h00;
RAM[16'h0B37] = 8'h00;
RAM[16'h0B38] = 8'h00;
RAM[16'h0B39] = 8'h00;
RAM[16'h0B3A] = 8'h00;
RAM[16'h0B3B] = 8'h00;
RAM[16'h0B3C] = 8'h00;
RAM[16'h0B3D] = 8'h00;
RAM[16'h0B3E] = 8'h00;
RAM[16'h0B3F] = 8'h00;
RAM[16'h0B40] = 8'h00;
RAM[16'h0B41] = 8'h00;
RAM[16'h0B42] = 8'h00;
RAM[16'h0B43] = 8'h00;
RAM[16'h0B44] = 8'h00;
RAM[16'h0B45] = 8'h00;
RAM[16'h0B46] = 8'h00;
RAM[16'h0B47] = 8'h00;
RAM[16'h0B48] = 8'h00;
RAM[16'h0B49] = 8'h00;
RAM[16'h0B4A] = 8'h00;
RAM[16'h0B4B] = 8'h00;
RAM[16'h0B4C] = 8'h00;
RAM[16'h0B4D] = 8'h00;
RAM[16'h0B4E] = 8'h00;
RAM[16'h0B4F] = 8'h00;
RAM[16'h0B50] = 8'h00;
RAM[16'h0B51] = 8'h00;
RAM[16'h0B52] = 8'h00;
RAM[16'h0B53] = 8'h00;
RAM[16'h0B54] = 8'h00;
RAM[16'h0B55] = 8'h00;
RAM[16'h0B56] = 8'h00;
RAM[16'h0B57] = 8'h00;
RAM[16'h0B58] = 8'h00;
RAM[16'h0B59] = 8'h00;
RAM[16'h0B5A] = 8'h00;
RAM[16'h0B5B] = 8'h00;
RAM[16'h0B5C] = 8'h00;
RAM[16'h0B5D] = 8'h00;
RAM[16'h0B5E] = 8'h00;
RAM[16'h0B5F] = 8'h00;
RAM[16'h0B60] = 8'h00;
RAM[16'h0B61] = 8'h00;
RAM[16'h0B62] = 8'h00;
RAM[16'h0B63] = 8'h00;
RAM[16'h0B64] = 8'h00;
RAM[16'h0B65] = 8'h00;
RAM[16'h0B66] = 8'h00;
RAM[16'h0B67] = 8'h00;
RAM[16'h0B68] = 8'h00;
RAM[16'h0B69] = 8'h00;
RAM[16'h0B6A] = 8'h00;
RAM[16'h0B6B] = 8'h00;
RAM[16'h0B6C] = 8'h00;
RAM[16'h0B6D] = 8'h00;
RAM[16'h0B6E] = 8'h00;
RAM[16'h0B6F] = 8'h00;
RAM[16'h0B70] = 8'h00;
RAM[16'h0B71] = 8'h00;
RAM[16'h0B72] = 8'h00;
RAM[16'h0B73] = 8'h00;
RAM[16'h0B74] = 8'h00;
RAM[16'h0B75] = 8'h00;
RAM[16'h0B76] = 8'h00;
RAM[16'h0B77] = 8'h00;
RAM[16'h0B78] = 8'h00;
RAM[16'h0B79] = 8'h00;
RAM[16'h0B7A] = 8'h00;
RAM[16'h0B7B] = 8'h00;
RAM[16'h0B7C] = 8'h00;
RAM[16'h0B7D] = 8'h00;
RAM[16'h0B7E] = 8'h00;
RAM[16'h0B7F] = 8'h00;
RAM[16'h0B80] = 8'h00;
RAM[16'h0B81] = 8'h00;
RAM[16'h0B82] = 8'h00;
RAM[16'h0B83] = 8'h00;
RAM[16'h0B84] = 8'h00;
RAM[16'h0B85] = 8'h00;
RAM[16'h0B86] = 8'h00;
RAM[16'h0B87] = 8'h00;
RAM[16'h0B88] = 8'h00;
RAM[16'h0B89] = 8'h00;
RAM[16'h0B8A] = 8'h00;
RAM[16'h0B8B] = 8'h00;
RAM[16'h0B8C] = 8'h00;
RAM[16'h0B8D] = 8'h00;
RAM[16'h0B8E] = 8'h00;
RAM[16'h0B8F] = 8'h00;
RAM[16'h0B90] = 8'h00;
RAM[16'h0B91] = 8'h00;
RAM[16'h0B92] = 8'h00;
RAM[16'h0B93] = 8'h00;
RAM[16'h0B94] = 8'h00;
RAM[16'h0B95] = 8'h00;
RAM[16'h0B96] = 8'h00;
RAM[16'h0B97] = 8'h00;
RAM[16'h0B98] = 8'h00;
RAM[16'h0B99] = 8'h00;
RAM[16'h0B9A] = 8'h00;
RAM[16'h0B9B] = 8'h00;
RAM[16'h0B9C] = 8'h00;
RAM[16'h0B9D] = 8'h00;
RAM[16'h0B9E] = 8'h00;
RAM[16'h0B9F] = 8'h00;
RAM[16'h0BA0] = 8'h00;
RAM[16'h0BA1] = 8'h00;
RAM[16'h0BA2] = 8'h00;
RAM[16'h0BA3] = 8'h00;
RAM[16'h0BA4] = 8'h00;
RAM[16'h0BA5] = 8'h00;
RAM[16'h0BA6] = 8'h00;
RAM[16'h0BA7] = 8'h00;
RAM[16'h0BA8] = 8'h00;
RAM[16'h0BA9] = 8'h00;
RAM[16'h0BAA] = 8'h00;
RAM[16'h0BAB] = 8'h00;
RAM[16'h0BAC] = 8'h00;
RAM[16'h0BAD] = 8'h00;
RAM[16'h0BAE] = 8'h00;
RAM[16'h0BAF] = 8'h00;
RAM[16'h0BB0] = 8'h00;
RAM[16'h0BB1] = 8'h00;
RAM[16'h0BB2] = 8'h00;
RAM[16'h0BB3] = 8'h00;
RAM[16'h0BB4] = 8'h00;
RAM[16'h0BB5] = 8'h00;
RAM[16'h0BB6] = 8'h00;
RAM[16'h0BB7] = 8'h00;
RAM[16'h0BB8] = 8'h00;
RAM[16'h0BB9] = 8'h00;
RAM[16'h0BBA] = 8'h00;
RAM[16'h0BBB] = 8'h00;
RAM[16'h0BBC] = 8'h00;
RAM[16'h0BBD] = 8'h00;
RAM[16'h0BBE] = 8'h00;
RAM[16'h0BBF] = 8'h00;
RAM[16'h0BC0] = 8'h00;
RAM[16'h0BC1] = 8'h00;
RAM[16'h0BC2] = 8'h00;
RAM[16'h0BC3] = 8'h00;
RAM[16'h0BC4] = 8'h00;
RAM[16'h0BC5] = 8'h00;
RAM[16'h0BC6] = 8'h00;
RAM[16'h0BC7] = 8'h00;
RAM[16'h0BC8] = 8'h00;
RAM[16'h0BC9] = 8'h00;
RAM[16'h0BCA] = 8'h00;
RAM[16'h0BCB] = 8'h00;
RAM[16'h0BCC] = 8'h00;
RAM[16'h0BCD] = 8'h00;
RAM[16'h0BCE] = 8'h00;
RAM[16'h0BCF] = 8'h00;
RAM[16'h0BD0] = 8'h00;
RAM[16'h0BD1] = 8'h00;
RAM[16'h0BD2] = 8'h00;
RAM[16'h0BD3] = 8'h00;
RAM[16'h0BD4] = 8'h00;
RAM[16'h0BD5] = 8'h00;
RAM[16'h0BD6] = 8'h00;
RAM[16'h0BD7] = 8'h00;
RAM[16'h0BD8] = 8'h00;
RAM[16'h0BD9] = 8'h00;
RAM[16'h0BDA] = 8'h00;
RAM[16'h0BDB] = 8'h00;
RAM[16'h0BDC] = 8'h00;
RAM[16'h0BDD] = 8'h00;
RAM[16'h0BDE] = 8'h00;
RAM[16'h0BDF] = 8'h00;
RAM[16'h0BE0] = 8'h00;
RAM[16'h0BE1] = 8'h00;
RAM[16'h0BE2] = 8'h00;
RAM[16'h0BE3] = 8'h00;
RAM[16'h0BE4] = 8'h00;
RAM[16'h0BE5] = 8'h00;
RAM[16'h0BE6] = 8'h00;
RAM[16'h0BE7] = 8'h00;
RAM[16'h0BE8] = 8'h00;
RAM[16'h0BE9] = 8'h00;
RAM[16'h0BEA] = 8'h00;
RAM[16'h0BEB] = 8'h00;
RAM[16'h0BEC] = 8'h00;
RAM[16'h0BED] = 8'h00;
RAM[16'h0BEE] = 8'h00;
RAM[16'h0BEF] = 8'h00;
RAM[16'h0BF0] = 8'h00;
RAM[16'h0BF1] = 8'h00;
RAM[16'h0BF2] = 8'h00;
RAM[16'h0BF3] = 8'h00;
RAM[16'h0BF4] = 8'h00;
RAM[16'h0BF5] = 8'h00;
RAM[16'h0BF6] = 8'h00;
RAM[16'h0BF7] = 8'h00;
RAM[16'h0BF8] = 8'h00;
RAM[16'h0BF9] = 8'h00;
RAM[16'h0BFA] = 8'h00;
RAM[16'h0BFB] = 8'h00;
RAM[16'h0BFC] = 8'h00;
RAM[16'h0BFD] = 8'h00;
RAM[16'h0BFE] = 8'h00;
RAM[16'h0BFF] = 8'h00;
RAM[16'h0C00] = 8'h00;
RAM[16'h0C01] = 8'h00;
RAM[16'h0C02] = 8'h00;
RAM[16'h0C03] = 8'h00;
RAM[16'h0C04] = 8'h00;
RAM[16'h0C05] = 8'h00;
RAM[16'h0C06] = 8'h00;
RAM[16'h0C07] = 8'h00;
RAM[16'h0C08] = 8'h00;
RAM[16'h0C09] = 8'h00;
RAM[16'h0C0A] = 8'h00;
RAM[16'h0C0B] = 8'h00;
RAM[16'h0C0C] = 8'h00;
RAM[16'h0C0D] = 8'h00;
RAM[16'h0C0E] = 8'h00;
RAM[16'h0C0F] = 8'h00;
RAM[16'h0C10] = 8'h00;
RAM[16'h0C11] = 8'h00;
RAM[16'h0C12] = 8'h00;
RAM[16'h0C13] = 8'h00;
RAM[16'h0C14] = 8'h00;
RAM[16'h0C15] = 8'h00;
RAM[16'h0C16] = 8'h00;
RAM[16'h0C17] = 8'h00;
RAM[16'h0C18] = 8'h00;
RAM[16'h0C19] = 8'h00;
RAM[16'h0C1A] = 8'h00;
RAM[16'h0C1B] = 8'h00;
RAM[16'h0C1C] = 8'h00;
RAM[16'h0C1D] = 8'h00;
RAM[16'h0C1E] = 8'h00;
RAM[16'h0C1F] = 8'h00;
RAM[16'h0C20] = 8'h00;
RAM[16'h0C21] = 8'h00;
RAM[16'h0C22] = 8'h00;
RAM[16'h0C23] = 8'h00;
RAM[16'h0C24] = 8'h00;
RAM[16'h0C25] = 8'h00;
RAM[16'h0C26] = 8'h00;
RAM[16'h0C27] = 8'h00;
RAM[16'h0C28] = 8'h00;
RAM[16'h0C29] = 8'h00;
RAM[16'h0C2A] = 8'h00;
RAM[16'h0C2B] = 8'h00;
RAM[16'h0C2C] = 8'h00;
RAM[16'h0C2D] = 8'h00;
RAM[16'h0C2E] = 8'h00;
RAM[16'h0C2F] = 8'h00;
RAM[16'h0C30] = 8'h00;
RAM[16'h0C31] = 8'h00;
RAM[16'h0C32] = 8'h00;
RAM[16'h0C33] = 8'h00;
RAM[16'h0C34] = 8'h00;
RAM[16'h0C35] = 8'h00;
RAM[16'h0C36] = 8'h00;
RAM[16'h0C37] = 8'h00;
RAM[16'h0C38] = 8'h00;
RAM[16'h0C39] = 8'h00;
RAM[16'h0C3A] = 8'h00;
RAM[16'h0C3B] = 8'h00;
RAM[16'h0C3C] = 8'h00;
RAM[16'h0C3D] = 8'h00;
RAM[16'h0C3E] = 8'h00;
RAM[16'h0C3F] = 8'h00;
RAM[16'h0C40] = 8'h00;
RAM[16'h0C41] = 8'h00;
RAM[16'h0C42] = 8'h00;
RAM[16'h0C43] = 8'h00;
RAM[16'h0C44] = 8'h00;
RAM[16'h0C45] = 8'h00;
RAM[16'h0C46] = 8'h00;
RAM[16'h0C47] = 8'h00;
RAM[16'h0C48] = 8'h00;
RAM[16'h0C49] = 8'h00;
RAM[16'h0C4A] = 8'h00;
RAM[16'h0C4B] = 8'h00;
RAM[16'h0C4C] = 8'h00;
RAM[16'h0C4D] = 8'h00;
RAM[16'h0C4E] = 8'h00;
RAM[16'h0C4F] = 8'h00;
RAM[16'h0C50] = 8'h00;
RAM[16'h0C51] = 8'h00;
RAM[16'h0C52] = 8'h00;
RAM[16'h0C53] = 8'h00;
RAM[16'h0C54] = 8'h00;
RAM[16'h0C55] = 8'h00;
RAM[16'h0C56] = 8'h00;
RAM[16'h0C57] = 8'h00;
RAM[16'h0C58] = 8'h00;
RAM[16'h0C59] = 8'h00;
RAM[16'h0C5A] = 8'h00;
RAM[16'h0C5B] = 8'h00;
RAM[16'h0C5C] = 8'h00;
RAM[16'h0C5D] = 8'h00;
RAM[16'h0C5E] = 8'h00;
RAM[16'h0C5F] = 8'h00;
RAM[16'h0C60] = 8'h00;
RAM[16'h0C61] = 8'h00;
RAM[16'h0C62] = 8'h00;
RAM[16'h0C63] = 8'h00;
RAM[16'h0C64] = 8'h00;
RAM[16'h0C65] = 8'h00;
RAM[16'h0C66] = 8'h00;
RAM[16'h0C67] = 8'h00;
RAM[16'h0C68] = 8'h00;
RAM[16'h0C69] = 8'h00;
RAM[16'h0C6A] = 8'h00;
RAM[16'h0C6B] = 8'h00;
RAM[16'h0C6C] = 8'h00;
RAM[16'h0C6D] = 8'h00;
RAM[16'h0C6E] = 8'h00;
RAM[16'h0C6F] = 8'h00;
RAM[16'h0C70] = 8'h00;
RAM[16'h0C71] = 8'h00;
RAM[16'h0C72] = 8'h00;
RAM[16'h0C73] = 8'h00;
RAM[16'h0C74] = 8'h00;
RAM[16'h0C75] = 8'h00;
RAM[16'h0C76] = 8'h00;
RAM[16'h0C77] = 8'h00;
RAM[16'h0C78] = 8'h00;
RAM[16'h0C79] = 8'h00;
RAM[16'h0C7A] = 8'h00;
RAM[16'h0C7B] = 8'h00;
RAM[16'h0C7C] = 8'h00;
RAM[16'h0C7D] = 8'h00;
RAM[16'h0C7E] = 8'h00;
RAM[16'h0C7F] = 8'h00;
RAM[16'h0C80] = 8'h00;
RAM[16'h0C81] = 8'h00;
RAM[16'h0C82] = 8'h00;
RAM[16'h0C83] = 8'h00;
RAM[16'h0C84] = 8'h00;
RAM[16'h0C85] = 8'h00;
RAM[16'h0C86] = 8'h00;
RAM[16'h0C87] = 8'h00;
RAM[16'h0C88] = 8'h00;
RAM[16'h0C89] = 8'h00;
RAM[16'h0C8A] = 8'h00;
RAM[16'h0C8B] = 8'h00;
RAM[16'h0C8C] = 8'h00;
RAM[16'h0C8D] = 8'h00;
RAM[16'h0C8E] = 8'h00;
RAM[16'h0C8F] = 8'h00;
RAM[16'h0C90] = 8'h00;
RAM[16'h0C91] = 8'h00;
RAM[16'h0C92] = 8'h00;
RAM[16'h0C93] = 8'h00;
RAM[16'h0C94] = 8'h00;
RAM[16'h0C95] = 8'h00;
RAM[16'h0C96] = 8'h00;
RAM[16'h0C97] = 8'h00;
RAM[16'h0C98] = 8'h00;
RAM[16'h0C99] = 8'h00;
RAM[16'h0C9A] = 8'h00;
RAM[16'h0C9B] = 8'h00;
RAM[16'h0C9C] = 8'h00;
RAM[16'h0C9D] = 8'h00;
RAM[16'h0C9E] = 8'h00;
RAM[16'h0C9F] = 8'h00;
RAM[16'h0CA0] = 8'h00;
RAM[16'h0CA1] = 8'h00;
RAM[16'h0CA2] = 8'h00;
RAM[16'h0CA3] = 8'h00;
RAM[16'h0CA4] = 8'h00;
RAM[16'h0CA5] = 8'h00;
RAM[16'h0CA6] = 8'h00;
RAM[16'h0CA7] = 8'h00;
RAM[16'h0CA8] = 8'h00;
RAM[16'h0CA9] = 8'h00;
RAM[16'h0CAA] = 8'h00;
RAM[16'h0CAB] = 8'h00;
RAM[16'h0CAC] = 8'h00;
RAM[16'h0CAD] = 8'h00;
RAM[16'h0CAE] = 8'h00;
RAM[16'h0CAF] = 8'h00;
RAM[16'h0CB0] = 8'h00;
RAM[16'h0CB1] = 8'h00;
RAM[16'h0CB2] = 8'h00;
RAM[16'h0CB3] = 8'h00;
RAM[16'h0CB4] = 8'h00;
RAM[16'h0CB5] = 8'h00;
RAM[16'h0CB6] = 8'h00;
RAM[16'h0CB7] = 8'h00;
RAM[16'h0CB8] = 8'h00;
RAM[16'h0CB9] = 8'h00;
RAM[16'h0CBA] = 8'h00;
RAM[16'h0CBB] = 8'h00;
RAM[16'h0CBC] = 8'h00;
RAM[16'h0CBD] = 8'h00;
RAM[16'h0CBE] = 8'h00;
RAM[16'h0CBF] = 8'h00;
RAM[16'h0CC0] = 8'h00;
RAM[16'h0CC1] = 8'h00;
RAM[16'h0CC2] = 8'h00;
RAM[16'h0CC3] = 8'h00;
RAM[16'h0CC4] = 8'h00;
RAM[16'h0CC5] = 8'h00;
RAM[16'h0CC6] = 8'h00;
RAM[16'h0CC7] = 8'h00;
RAM[16'h0CC8] = 8'h00;
RAM[16'h0CC9] = 8'h00;
RAM[16'h0CCA] = 8'h00;
RAM[16'h0CCB] = 8'h00;
RAM[16'h0CCC] = 8'h00;
RAM[16'h0CCD] = 8'h00;
RAM[16'h0CCE] = 8'h00;
RAM[16'h0CCF] = 8'h00;
RAM[16'h0CD0] = 8'h00;
RAM[16'h0CD1] = 8'h00;
RAM[16'h0CD2] = 8'h00;
RAM[16'h0CD3] = 8'h00;
RAM[16'h0CD4] = 8'h00;
RAM[16'h0CD5] = 8'h00;
RAM[16'h0CD6] = 8'h00;
RAM[16'h0CD7] = 8'h00;
RAM[16'h0CD8] = 8'h00;
RAM[16'h0CD9] = 8'h00;
RAM[16'h0CDA] = 8'h00;
RAM[16'h0CDB] = 8'h00;
RAM[16'h0CDC] = 8'h00;
RAM[16'h0CDD] = 8'h00;
RAM[16'h0CDE] = 8'h00;
RAM[16'h0CDF] = 8'h00;
RAM[16'h0CE0] = 8'h00;
RAM[16'h0CE1] = 8'h00;
RAM[16'h0CE2] = 8'h00;
RAM[16'h0CE3] = 8'h00;
RAM[16'h0CE4] = 8'h00;
RAM[16'h0CE5] = 8'h00;
RAM[16'h0CE6] = 8'h00;
RAM[16'h0CE7] = 8'h00;
RAM[16'h0CE8] = 8'h00;
RAM[16'h0CE9] = 8'h00;
RAM[16'h0CEA] = 8'h00;
RAM[16'h0CEB] = 8'h00;
RAM[16'h0CEC] = 8'h00;
RAM[16'h0CED] = 8'h00;
RAM[16'h0CEE] = 8'h00;
RAM[16'h0CEF] = 8'h00;
RAM[16'h0CF0] = 8'h00;
RAM[16'h0CF1] = 8'h00;
RAM[16'h0CF2] = 8'h00;
RAM[16'h0CF3] = 8'h00;
RAM[16'h0CF4] = 8'h00;
RAM[16'h0CF5] = 8'h00;
RAM[16'h0CF6] = 8'h00;
RAM[16'h0CF7] = 8'h00;
RAM[16'h0CF8] = 8'h00;
RAM[16'h0CF9] = 8'h00;
RAM[16'h0CFA] = 8'h00;
RAM[16'h0CFB] = 8'h00;
RAM[16'h0CFC] = 8'h00;
RAM[16'h0CFD] = 8'h00;
RAM[16'h0CFE] = 8'h00;
RAM[16'h0CFF] = 8'h00;
RAM[16'h0D00] = 8'h00;
RAM[16'h0D01] = 8'h00;
RAM[16'h0D02] = 8'h00;
RAM[16'h0D03] = 8'h00;
RAM[16'h0D04] = 8'h00;
RAM[16'h0D05] = 8'h00;
RAM[16'h0D06] = 8'h00;
RAM[16'h0D07] = 8'h00;
RAM[16'h0D08] = 8'h00;
RAM[16'h0D09] = 8'h00;
RAM[16'h0D0A] = 8'h00;
RAM[16'h0D0B] = 8'h00;
RAM[16'h0D0C] = 8'h00;
RAM[16'h0D0D] = 8'h00;
RAM[16'h0D0E] = 8'h00;
RAM[16'h0D0F] = 8'h00;
RAM[16'h0D10] = 8'h00;
RAM[16'h0D11] = 8'h00;
RAM[16'h0D12] = 8'h00;
RAM[16'h0D13] = 8'h00;
RAM[16'h0D14] = 8'h00;
RAM[16'h0D15] = 8'h00;
RAM[16'h0D16] = 8'h00;
RAM[16'h0D17] = 8'h00;
RAM[16'h0D18] = 8'h00;
RAM[16'h0D19] = 8'h00;
RAM[16'h0D1A] = 8'h00;
RAM[16'h0D1B] = 8'h00;
RAM[16'h0D1C] = 8'h00;
RAM[16'h0D1D] = 8'h00;
RAM[16'h0D1E] = 8'h00;
RAM[16'h0D1F] = 8'h00;
RAM[16'h0D20] = 8'h00;
RAM[16'h0D21] = 8'h00;
RAM[16'h0D22] = 8'h00;
RAM[16'h0D23] = 8'h00;
RAM[16'h0D24] = 8'h00;
RAM[16'h0D25] = 8'h00;
RAM[16'h0D26] = 8'h00;
RAM[16'h0D27] = 8'h00;
RAM[16'h0D28] = 8'h00;
RAM[16'h0D29] = 8'h00;
RAM[16'h0D2A] = 8'h00;
RAM[16'h0D2B] = 8'h00;
RAM[16'h0D2C] = 8'h00;
RAM[16'h0D2D] = 8'h00;
RAM[16'h0D2E] = 8'h00;
RAM[16'h0D2F] = 8'h00;
RAM[16'h0D30] = 8'h00;
RAM[16'h0D31] = 8'h00;
RAM[16'h0D32] = 8'h00;
RAM[16'h0D33] = 8'h00;
RAM[16'h0D34] = 8'h00;
RAM[16'h0D35] = 8'h00;
RAM[16'h0D36] = 8'h00;
RAM[16'h0D37] = 8'h00;
RAM[16'h0D38] = 8'h00;
RAM[16'h0D39] = 8'h00;
RAM[16'h0D3A] = 8'h00;
RAM[16'h0D3B] = 8'h00;
RAM[16'h0D3C] = 8'h00;
RAM[16'h0D3D] = 8'h00;
RAM[16'h0D3E] = 8'h00;
RAM[16'h0D3F] = 8'h00;
RAM[16'h0D40] = 8'h00;
RAM[16'h0D41] = 8'h00;
RAM[16'h0D42] = 8'h00;
RAM[16'h0D43] = 8'h00;
RAM[16'h0D44] = 8'h00;
RAM[16'h0D45] = 8'h00;
RAM[16'h0D46] = 8'h00;
RAM[16'h0D47] = 8'h00;
RAM[16'h0D48] = 8'h00;
RAM[16'h0D49] = 8'h00;
RAM[16'h0D4A] = 8'h00;
RAM[16'h0D4B] = 8'h00;
RAM[16'h0D4C] = 8'h00;
RAM[16'h0D4D] = 8'h00;
RAM[16'h0D4E] = 8'h00;
RAM[16'h0D4F] = 8'h00;
RAM[16'h0D50] = 8'h00;
RAM[16'h0D51] = 8'h00;
RAM[16'h0D52] = 8'h00;
RAM[16'h0D53] = 8'h00;
RAM[16'h0D54] = 8'h00;
RAM[16'h0D55] = 8'h00;
RAM[16'h0D56] = 8'h00;
RAM[16'h0D57] = 8'h00;
RAM[16'h0D58] = 8'h00;
RAM[16'h0D59] = 8'h00;
RAM[16'h0D5A] = 8'h00;
RAM[16'h0D5B] = 8'h00;
RAM[16'h0D5C] = 8'h00;
RAM[16'h0D5D] = 8'h00;
RAM[16'h0D5E] = 8'h00;
RAM[16'h0D5F] = 8'h00;
RAM[16'h0D60] = 8'h00;
RAM[16'h0D61] = 8'h00;
RAM[16'h0D62] = 8'h00;
RAM[16'h0D63] = 8'h00;
RAM[16'h0D64] = 8'h00;
RAM[16'h0D65] = 8'h00;
RAM[16'h0D66] = 8'h00;
RAM[16'h0D67] = 8'h00;
RAM[16'h0D68] = 8'h00;
RAM[16'h0D69] = 8'h00;
RAM[16'h0D6A] = 8'h00;
RAM[16'h0D6B] = 8'h00;
RAM[16'h0D6C] = 8'h00;
RAM[16'h0D6D] = 8'h00;
RAM[16'h0D6E] = 8'h00;
RAM[16'h0D6F] = 8'h00;
RAM[16'h0D70] = 8'h00;
RAM[16'h0D71] = 8'h00;
RAM[16'h0D72] = 8'h00;
RAM[16'h0D73] = 8'h00;
RAM[16'h0D74] = 8'h00;
RAM[16'h0D75] = 8'h00;
RAM[16'h0D76] = 8'h00;
RAM[16'h0D77] = 8'h00;
RAM[16'h0D78] = 8'h00;
RAM[16'h0D79] = 8'h00;
RAM[16'h0D7A] = 8'h00;
RAM[16'h0D7B] = 8'h00;
RAM[16'h0D7C] = 8'h00;
RAM[16'h0D7D] = 8'h00;
RAM[16'h0D7E] = 8'h00;
RAM[16'h0D7F] = 8'h00;
RAM[16'h0D80] = 8'h00;
RAM[16'h0D81] = 8'h00;
RAM[16'h0D82] = 8'h00;
RAM[16'h0D83] = 8'h00;
RAM[16'h0D84] = 8'h00;
RAM[16'h0D85] = 8'h00;
RAM[16'h0D86] = 8'h00;
RAM[16'h0D87] = 8'h00;
RAM[16'h0D88] = 8'h00;
RAM[16'h0D89] = 8'h00;
RAM[16'h0D8A] = 8'h00;
RAM[16'h0D8B] = 8'h00;
RAM[16'h0D8C] = 8'h00;
RAM[16'h0D8D] = 8'h00;
RAM[16'h0D8E] = 8'h00;
RAM[16'h0D8F] = 8'h00;
RAM[16'h0D90] = 8'h00;
RAM[16'h0D91] = 8'h00;
RAM[16'h0D92] = 8'h00;
RAM[16'h0D93] = 8'h00;
RAM[16'h0D94] = 8'h00;
RAM[16'h0D95] = 8'h00;
RAM[16'h0D96] = 8'h00;
RAM[16'h0D97] = 8'h00;
RAM[16'h0D98] = 8'h00;
RAM[16'h0D99] = 8'h00;
RAM[16'h0D9A] = 8'h00;
RAM[16'h0D9B] = 8'h00;
RAM[16'h0D9C] = 8'h00;
RAM[16'h0D9D] = 8'h00;
RAM[16'h0D9E] = 8'h00;
RAM[16'h0D9F] = 8'h00;
RAM[16'h0DA0] = 8'h00;
RAM[16'h0DA1] = 8'h00;
RAM[16'h0DA2] = 8'h00;
RAM[16'h0DA3] = 8'h00;
RAM[16'h0DA4] = 8'h00;
RAM[16'h0DA5] = 8'h00;
RAM[16'h0DA6] = 8'h00;
RAM[16'h0DA7] = 8'h00;
RAM[16'h0DA8] = 8'h00;
RAM[16'h0DA9] = 8'h00;
RAM[16'h0DAA] = 8'h00;
RAM[16'h0DAB] = 8'h00;
RAM[16'h0DAC] = 8'h00;
RAM[16'h0DAD] = 8'h00;
RAM[16'h0DAE] = 8'h00;
RAM[16'h0DAF] = 8'h00;
RAM[16'h0DB0] = 8'h00;
RAM[16'h0DB1] = 8'h00;
RAM[16'h0DB2] = 8'h00;
RAM[16'h0DB3] = 8'h00;
RAM[16'h0DB4] = 8'h00;
RAM[16'h0DB5] = 8'h00;
RAM[16'h0DB6] = 8'h00;
RAM[16'h0DB7] = 8'h00;
RAM[16'h0DB8] = 8'h00;
RAM[16'h0DB9] = 8'h00;
RAM[16'h0DBA] = 8'h00;
RAM[16'h0DBB] = 8'h00;
RAM[16'h0DBC] = 8'h00;
RAM[16'h0DBD] = 8'h00;
RAM[16'h0DBE] = 8'h00;
RAM[16'h0DBF] = 8'h00;
RAM[16'h0DC0] = 8'h00;
RAM[16'h0DC1] = 8'h00;
RAM[16'h0DC2] = 8'h00;
RAM[16'h0DC3] = 8'h00;
RAM[16'h0DC4] = 8'h00;
RAM[16'h0DC5] = 8'h00;
RAM[16'h0DC6] = 8'h00;
RAM[16'h0DC7] = 8'h00;
RAM[16'h0DC8] = 8'h00;
RAM[16'h0DC9] = 8'h00;
RAM[16'h0DCA] = 8'h00;
RAM[16'h0DCB] = 8'h00;
RAM[16'h0DCC] = 8'h00;
RAM[16'h0DCD] = 8'h00;
RAM[16'h0DCE] = 8'h00;
RAM[16'h0DCF] = 8'h00;
RAM[16'h0DD0] = 8'h00;
RAM[16'h0DD1] = 8'h00;
RAM[16'h0DD2] = 8'h00;
RAM[16'h0DD3] = 8'h00;
RAM[16'h0DD4] = 8'h00;
RAM[16'h0DD5] = 8'h00;
RAM[16'h0DD6] = 8'h00;
RAM[16'h0DD7] = 8'h00;
RAM[16'h0DD8] = 8'h00;
RAM[16'h0DD9] = 8'h00;
RAM[16'h0DDA] = 8'h00;
RAM[16'h0DDB] = 8'h00;
RAM[16'h0DDC] = 8'h00;
RAM[16'h0DDD] = 8'h00;
RAM[16'h0DDE] = 8'h00;
RAM[16'h0DDF] = 8'h00;
RAM[16'h0DE0] = 8'h00;
RAM[16'h0DE1] = 8'h00;
RAM[16'h0DE2] = 8'h00;
RAM[16'h0DE3] = 8'h00;
RAM[16'h0DE4] = 8'h00;
RAM[16'h0DE5] = 8'h00;
RAM[16'h0DE6] = 8'h00;
RAM[16'h0DE7] = 8'h00;
RAM[16'h0DE8] = 8'h00;
RAM[16'h0DE9] = 8'h00;
RAM[16'h0DEA] = 8'h00;
RAM[16'h0DEB] = 8'h00;
RAM[16'h0DEC] = 8'h00;
RAM[16'h0DED] = 8'h00;
RAM[16'h0DEE] = 8'h00;
RAM[16'h0DEF] = 8'h00;
RAM[16'h0DF0] = 8'h00;
RAM[16'h0DF1] = 8'h00;
RAM[16'h0DF2] = 8'h00;
RAM[16'h0DF3] = 8'h00;
RAM[16'h0DF4] = 8'h00;
RAM[16'h0DF5] = 8'h00;
RAM[16'h0DF6] = 8'h00;
RAM[16'h0DF7] = 8'h00;
RAM[16'h0DF8] = 8'h00;
RAM[16'h0DF9] = 8'h00;
RAM[16'h0DFA] = 8'h00;
RAM[16'h0DFB] = 8'h00;
RAM[16'h0DFC] = 8'h00;
RAM[16'h0DFD] = 8'h00;
RAM[16'h0DFE] = 8'h00;
RAM[16'h0DFF] = 8'h00;
RAM[16'h0E00] = 8'h00;
RAM[16'h0E01] = 8'h00;
RAM[16'h0E02] = 8'h00;
RAM[16'h0E03] = 8'h00;
RAM[16'h0E04] = 8'h00;
RAM[16'h0E05] = 8'h00;
RAM[16'h0E06] = 8'h00;
RAM[16'h0E07] = 8'h00;
RAM[16'h0E08] = 8'h00;
RAM[16'h0E09] = 8'h00;
RAM[16'h0E0A] = 8'h00;
RAM[16'h0E0B] = 8'h00;
RAM[16'h0E0C] = 8'h00;
RAM[16'h0E0D] = 8'h00;
RAM[16'h0E0E] = 8'h00;
RAM[16'h0E0F] = 8'h00;
RAM[16'h0E10] = 8'h00;
RAM[16'h0E11] = 8'h00;
RAM[16'h0E12] = 8'h00;
RAM[16'h0E13] = 8'h00;
RAM[16'h0E14] = 8'h00;
RAM[16'h0E15] = 8'h00;
RAM[16'h0E16] = 8'h00;
RAM[16'h0E17] = 8'h00;
RAM[16'h0E18] = 8'h00;
RAM[16'h0E19] = 8'h00;
RAM[16'h0E1A] = 8'h00;
RAM[16'h0E1B] = 8'h00;
RAM[16'h0E1C] = 8'h00;
RAM[16'h0E1D] = 8'h00;
RAM[16'h0E1E] = 8'h00;
RAM[16'h0E1F] = 8'h00;
RAM[16'h0E20] = 8'h00;
RAM[16'h0E21] = 8'h00;
RAM[16'h0E22] = 8'h00;
RAM[16'h0E23] = 8'h00;
RAM[16'h0E24] = 8'h00;
RAM[16'h0E25] = 8'h00;
RAM[16'h0E26] = 8'h00;
RAM[16'h0E27] = 8'h00;
RAM[16'h0E28] = 8'h00;
RAM[16'h0E29] = 8'h00;
RAM[16'h0E2A] = 8'h00;
RAM[16'h0E2B] = 8'h00;
RAM[16'h0E2C] = 8'h00;
RAM[16'h0E2D] = 8'h00;
RAM[16'h0E2E] = 8'h00;
RAM[16'h0E2F] = 8'h00;
RAM[16'h0E30] = 8'h00;
RAM[16'h0E31] = 8'h00;
RAM[16'h0E32] = 8'h00;
RAM[16'h0E33] = 8'h00;
RAM[16'h0E34] = 8'h00;
RAM[16'h0E35] = 8'h00;
RAM[16'h0E36] = 8'h00;
RAM[16'h0E37] = 8'h00;
RAM[16'h0E38] = 8'h00;
RAM[16'h0E39] = 8'h00;
RAM[16'h0E3A] = 8'h00;
RAM[16'h0E3B] = 8'h00;
RAM[16'h0E3C] = 8'h00;
RAM[16'h0E3D] = 8'h00;
RAM[16'h0E3E] = 8'h00;
RAM[16'h0E3F] = 8'h00;
RAM[16'h0E40] = 8'h00;
RAM[16'h0E41] = 8'h00;
RAM[16'h0E42] = 8'h00;
RAM[16'h0E43] = 8'h00;
RAM[16'h0E44] = 8'h00;
RAM[16'h0E45] = 8'h00;
RAM[16'h0E46] = 8'h00;
RAM[16'h0E47] = 8'h00;
RAM[16'h0E48] = 8'h00;
RAM[16'h0E49] = 8'h00;
RAM[16'h0E4A] = 8'h00;
RAM[16'h0E4B] = 8'h00;
RAM[16'h0E4C] = 8'h00;
RAM[16'h0E4D] = 8'h00;
RAM[16'h0E4E] = 8'h00;
RAM[16'h0E4F] = 8'h00;
RAM[16'h0E50] = 8'h00;
RAM[16'h0E51] = 8'h00;
RAM[16'h0E52] = 8'h00;
RAM[16'h0E53] = 8'h00;
RAM[16'h0E54] = 8'h00;
RAM[16'h0E55] = 8'h00;
RAM[16'h0E56] = 8'h00;
RAM[16'h0E57] = 8'h00;
RAM[16'h0E58] = 8'h00;
RAM[16'h0E59] = 8'h00;
RAM[16'h0E5A] = 8'h00;
RAM[16'h0E5B] = 8'h00;
RAM[16'h0E5C] = 8'h00;
RAM[16'h0E5D] = 8'h00;
RAM[16'h0E5E] = 8'h00;
RAM[16'h0E5F] = 8'h00;
RAM[16'h0E60] = 8'h00;
RAM[16'h0E61] = 8'h00;
RAM[16'h0E62] = 8'h00;
RAM[16'h0E63] = 8'h00;
RAM[16'h0E64] = 8'h00;
RAM[16'h0E65] = 8'h00;
RAM[16'h0E66] = 8'h00;
RAM[16'h0E67] = 8'h00;
RAM[16'h0E68] = 8'h00;
RAM[16'h0E69] = 8'h00;
RAM[16'h0E6A] = 8'h00;
RAM[16'h0E6B] = 8'h00;
RAM[16'h0E6C] = 8'h00;
RAM[16'h0E6D] = 8'h00;
RAM[16'h0E6E] = 8'h00;
RAM[16'h0E6F] = 8'h00;
RAM[16'h0E70] = 8'h00;
RAM[16'h0E71] = 8'h00;
RAM[16'h0E72] = 8'h00;
RAM[16'h0E73] = 8'h00;
RAM[16'h0E74] = 8'h00;
RAM[16'h0E75] = 8'h00;
RAM[16'h0E76] = 8'h00;
RAM[16'h0E77] = 8'h00;
RAM[16'h0E78] = 8'h00;
RAM[16'h0E79] = 8'h00;
RAM[16'h0E7A] = 8'h00;
RAM[16'h0E7B] = 8'h00;
RAM[16'h0E7C] = 8'h00;
RAM[16'h0E7D] = 8'h00;
RAM[16'h0E7E] = 8'h00;
RAM[16'h0E7F] = 8'h00;
RAM[16'h0E80] = 8'h00;
RAM[16'h0E81] = 8'h00;
RAM[16'h0E82] = 8'h00;
RAM[16'h0E83] = 8'h00;
RAM[16'h0E84] = 8'h00;
RAM[16'h0E85] = 8'h00;
RAM[16'h0E86] = 8'h00;
RAM[16'h0E87] = 8'h00;
RAM[16'h0E88] = 8'h00;
RAM[16'h0E89] = 8'h00;
RAM[16'h0E8A] = 8'h00;
RAM[16'h0E8B] = 8'h00;
RAM[16'h0E8C] = 8'h00;
RAM[16'h0E8D] = 8'h00;
RAM[16'h0E8E] = 8'h00;
RAM[16'h0E8F] = 8'h00;
RAM[16'h0E90] = 8'h00;
RAM[16'h0E91] = 8'h00;
RAM[16'h0E92] = 8'h00;
RAM[16'h0E93] = 8'h00;
RAM[16'h0E94] = 8'h00;
RAM[16'h0E95] = 8'h00;
RAM[16'h0E96] = 8'h00;
RAM[16'h0E97] = 8'h00;
RAM[16'h0E98] = 8'h00;
RAM[16'h0E99] = 8'h00;
RAM[16'h0E9A] = 8'h00;
RAM[16'h0E9B] = 8'h00;
RAM[16'h0E9C] = 8'h00;
RAM[16'h0E9D] = 8'h00;
RAM[16'h0E9E] = 8'h00;
RAM[16'h0E9F] = 8'h00;
RAM[16'h0EA0] = 8'h00;
RAM[16'h0EA1] = 8'h00;
RAM[16'h0EA2] = 8'h00;
RAM[16'h0EA3] = 8'h00;
RAM[16'h0EA4] = 8'h00;
RAM[16'h0EA5] = 8'h00;
RAM[16'h0EA6] = 8'h00;
RAM[16'h0EA7] = 8'h00;
RAM[16'h0EA8] = 8'h00;
RAM[16'h0EA9] = 8'h00;
RAM[16'h0EAA] = 8'h00;
RAM[16'h0EAB] = 8'h00;
RAM[16'h0EAC] = 8'h00;
RAM[16'h0EAD] = 8'h00;
RAM[16'h0EAE] = 8'h00;
RAM[16'h0EAF] = 8'h00;
RAM[16'h0EB0] = 8'h00;
RAM[16'h0EB1] = 8'h00;
RAM[16'h0EB2] = 8'h00;
RAM[16'h0EB3] = 8'h00;
RAM[16'h0EB4] = 8'h00;
RAM[16'h0EB5] = 8'h00;
RAM[16'h0EB6] = 8'h00;
RAM[16'h0EB7] = 8'h00;
RAM[16'h0EB8] = 8'h00;
RAM[16'h0EB9] = 8'h00;
RAM[16'h0EBA] = 8'h00;
RAM[16'h0EBB] = 8'h00;
RAM[16'h0EBC] = 8'h00;
RAM[16'h0EBD] = 8'h00;
RAM[16'h0EBE] = 8'h00;
RAM[16'h0EBF] = 8'h00;
RAM[16'h0EC0] = 8'h00;
RAM[16'h0EC1] = 8'h00;
RAM[16'h0EC2] = 8'h00;
RAM[16'h0EC3] = 8'h00;
RAM[16'h0EC4] = 8'h00;
RAM[16'h0EC5] = 8'h00;
RAM[16'h0EC6] = 8'h00;
RAM[16'h0EC7] = 8'h00;
RAM[16'h0EC8] = 8'h00;
RAM[16'h0EC9] = 8'h00;
RAM[16'h0ECA] = 8'h00;
RAM[16'h0ECB] = 8'h00;
RAM[16'h0ECC] = 8'h00;
RAM[16'h0ECD] = 8'h00;
RAM[16'h0ECE] = 8'h00;
RAM[16'h0ECF] = 8'h00;
RAM[16'h0ED0] = 8'h00;
RAM[16'h0ED1] = 8'h00;
RAM[16'h0ED2] = 8'h00;
RAM[16'h0ED3] = 8'h00;
RAM[16'h0ED4] = 8'h00;
RAM[16'h0ED5] = 8'h00;
RAM[16'h0ED6] = 8'h00;
RAM[16'h0ED7] = 8'h00;
RAM[16'h0ED8] = 8'h00;
RAM[16'h0ED9] = 8'h00;
RAM[16'h0EDA] = 8'h00;
RAM[16'h0EDB] = 8'h00;
RAM[16'h0EDC] = 8'h00;
RAM[16'h0EDD] = 8'h00;
RAM[16'h0EDE] = 8'h00;
RAM[16'h0EDF] = 8'h00;
RAM[16'h0EE0] = 8'h00;
RAM[16'h0EE1] = 8'h00;
RAM[16'h0EE2] = 8'h00;
RAM[16'h0EE3] = 8'h00;
RAM[16'h0EE4] = 8'h00;
RAM[16'h0EE5] = 8'h00;
RAM[16'h0EE6] = 8'h00;
RAM[16'h0EE7] = 8'h00;
RAM[16'h0EE8] = 8'h00;
RAM[16'h0EE9] = 8'h00;
RAM[16'h0EEA] = 8'h00;
RAM[16'h0EEB] = 8'h00;
RAM[16'h0EEC] = 8'h00;
RAM[16'h0EED] = 8'h00;
RAM[16'h0EEE] = 8'h00;
RAM[16'h0EEF] = 8'h00;
RAM[16'h0EF0] = 8'h00;
RAM[16'h0EF1] = 8'h00;
RAM[16'h0EF2] = 8'h00;
RAM[16'h0EF3] = 8'h00;
RAM[16'h0EF4] = 8'h00;
RAM[16'h0EF5] = 8'h00;
RAM[16'h0EF6] = 8'h00;
RAM[16'h0EF7] = 8'h00;
RAM[16'h0EF8] = 8'h00;
RAM[16'h0EF9] = 8'h00;
RAM[16'h0EFA] = 8'h00;
RAM[16'h0EFB] = 8'h00;
RAM[16'h0EFC] = 8'h00;
RAM[16'h0EFD] = 8'h00;
RAM[16'h0EFE] = 8'h00;
RAM[16'h0EFF] = 8'h00;
RAM[16'h0F00] = 8'h00;
RAM[16'h0F01] = 8'h00;
RAM[16'h0F02] = 8'h00;
RAM[16'h0F03] = 8'h00;
RAM[16'h0F04] = 8'h00;
RAM[16'h0F05] = 8'h00;
RAM[16'h0F06] = 8'h00;
RAM[16'h0F07] = 8'h00;
RAM[16'h0F08] = 8'h00;
RAM[16'h0F09] = 8'h00;
RAM[16'h0F0A] = 8'h00;
RAM[16'h0F0B] = 8'h00;
RAM[16'h0F0C] = 8'h00;
RAM[16'h0F0D] = 8'h00;
RAM[16'h0F0E] = 8'h00;
RAM[16'h0F0F] = 8'h00;
RAM[16'h0F10] = 8'h00;
RAM[16'h0F11] = 8'h00;
RAM[16'h0F12] = 8'h00;
RAM[16'h0F13] = 8'h00;
RAM[16'h0F14] = 8'h00;
RAM[16'h0F15] = 8'h00;
RAM[16'h0F16] = 8'h00;
RAM[16'h0F17] = 8'h00;
RAM[16'h0F18] = 8'h00;
RAM[16'h0F19] = 8'h00;
RAM[16'h0F1A] = 8'h00;
RAM[16'h0F1B] = 8'h00;
RAM[16'h0F1C] = 8'h00;
RAM[16'h0F1D] = 8'h00;
RAM[16'h0F1E] = 8'h00;
RAM[16'h0F1F] = 8'h00;
RAM[16'h0F20] = 8'h00;
RAM[16'h0F21] = 8'h00;
RAM[16'h0F22] = 8'h00;
RAM[16'h0F23] = 8'h00;
RAM[16'h0F24] = 8'h00;
RAM[16'h0F25] = 8'h00;
RAM[16'h0F26] = 8'h00;
RAM[16'h0F27] = 8'h00;
RAM[16'h0F28] = 8'h00;
RAM[16'h0F29] = 8'h00;
RAM[16'h0F2A] = 8'h00;
RAM[16'h0F2B] = 8'h00;
RAM[16'h0F2C] = 8'h00;
RAM[16'h0F2D] = 8'h00;
RAM[16'h0F2E] = 8'h00;
RAM[16'h0F2F] = 8'h00;
RAM[16'h0F30] = 8'h00;
RAM[16'h0F31] = 8'h00;
RAM[16'h0F32] = 8'h00;
RAM[16'h0F33] = 8'h00;
RAM[16'h0F34] = 8'h00;
RAM[16'h0F35] = 8'h00;
RAM[16'h0F36] = 8'h00;
RAM[16'h0F37] = 8'h00;
RAM[16'h0F38] = 8'h00;
RAM[16'h0F39] = 8'h00;
RAM[16'h0F3A] = 8'h00;
RAM[16'h0F3B] = 8'h00;
RAM[16'h0F3C] = 8'h00;
RAM[16'h0F3D] = 8'h00;
RAM[16'h0F3E] = 8'h00;
RAM[16'h0F3F] = 8'h00;
RAM[16'h0F40] = 8'h00;
RAM[16'h0F41] = 8'h00;
RAM[16'h0F42] = 8'h00;
RAM[16'h0F43] = 8'h00;
RAM[16'h0F44] = 8'h00;
RAM[16'h0F45] = 8'h00;
RAM[16'h0F46] = 8'h00;
RAM[16'h0F47] = 8'h00;
RAM[16'h0F48] = 8'h00;
RAM[16'h0F49] = 8'h00;
RAM[16'h0F4A] = 8'h00;
RAM[16'h0F4B] = 8'h00;
RAM[16'h0F4C] = 8'h00;
RAM[16'h0F4D] = 8'h00;
RAM[16'h0F4E] = 8'h00;
RAM[16'h0F4F] = 8'h00;
RAM[16'h0F50] = 8'h00;
RAM[16'h0F51] = 8'h00;
RAM[16'h0F52] = 8'h00;
RAM[16'h0F53] = 8'h00;
RAM[16'h0F54] = 8'h00;
RAM[16'h0F55] = 8'h00;
RAM[16'h0F56] = 8'h00;
RAM[16'h0F57] = 8'h00;
RAM[16'h0F58] = 8'h00;
RAM[16'h0F59] = 8'h00;
RAM[16'h0F5A] = 8'h00;
RAM[16'h0F5B] = 8'h00;
RAM[16'h0F5C] = 8'h00;
RAM[16'h0F5D] = 8'h00;
RAM[16'h0F5E] = 8'h00;
RAM[16'h0F5F] = 8'h00;
RAM[16'h0F60] = 8'h00;
RAM[16'h0F61] = 8'h00;
RAM[16'h0F62] = 8'h00;
RAM[16'h0F63] = 8'h00;
RAM[16'h0F64] = 8'h00;
RAM[16'h0F65] = 8'h00;
RAM[16'h0F66] = 8'h00;
RAM[16'h0F67] = 8'h00;
RAM[16'h0F68] = 8'h00;
RAM[16'h0F69] = 8'h00;
RAM[16'h0F6A] = 8'h00;
RAM[16'h0F6B] = 8'h00;
RAM[16'h0F6C] = 8'h00;
RAM[16'h0F6D] = 8'h00;
RAM[16'h0F6E] = 8'h00;
RAM[16'h0F6F] = 8'h00;
RAM[16'h0F70] = 8'h00;
RAM[16'h0F71] = 8'h00;
RAM[16'h0F72] = 8'h00;
RAM[16'h0F73] = 8'h00;
RAM[16'h0F74] = 8'h00;
RAM[16'h0F75] = 8'h00;
RAM[16'h0F76] = 8'h00;
RAM[16'h0F77] = 8'h00;
RAM[16'h0F78] = 8'h00;
RAM[16'h0F79] = 8'h00;
RAM[16'h0F7A] = 8'h00;
RAM[16'h0F7B] = 8'h00;
RAM[16'h0F7C] = 8'h00;
RAM[16'h0F7D] = 8'h00;
RAM[16'h0F7E] = 8'h00;
RAM[16'h0F7F] = 8'h00;
RAM[16'h0F80] = 8'h00;
RAM[16'h0F81] = 8'h00;
RAM[16'h0F82] = 8'h00;
RAM[16'h0F83] = 8'h00;
RAM[16'h0F84] = 8'h00;
RAM[16'h0F85] = 8'h00;
RAM[16'h0F86] = 8'h00;
RAM[16'h0F87] = 8'h00;
RAM[16'h0F88] = 8'h00;
RAM[16'h0F89] = 8'h00;
RAM[16'h0F8A] = 8'h00;
RAM[16'h0F8B] = 8'h00;
RAM[16'h0F8C] = 8'h00;
RAM[16'h0F8D] = 8'h00;
RAM[16'h0F8E] = 8'h00;
RAM[16'h0F8F] = 8'h00;
RAM[16'h0F90] = 8'h00;
RAM[16'h0F91] = 8'h00;
RAM[16'h0F92] = 8'h00;
RAM[16'h0F93] = 8'h00;
RAM[16'h0F94] = 8'h00;
RAM[16'h0F95] = 8'h00;
RAM[16'h0F96] = 8'h00;
RAM[16'h0F97] = 8'h00;
RAM[16'h0F98] = 8'h00;
RAM[16'h0F99] = 8'h00;
RAM[16'h0F9A] = 8'h00;
RAM[16'h0F9B] = 8'h00;
RAM[16'h0F9C] = 8'h00;
RAM[16'h0F9D] = 8'h00;
RAM[16'h0F9E] = 8'h00;
RAM[16'h0F9F] = 8'h00;
RAM[16'h0FA0] = 8'h00;
RAM[16'h0FA1] = 8'h00;
RAM[16'h0FA2] = 8'h00;
RAM[16'h0FA3] = 8'h00;
RAM[16'h0FA4] = 8'h00;
RAM[16'h0FA5] = 8'h00;
RAM[16'h0FA6] = 8'h00;
RAM[16'h0FA7] = 8'h00;
RAM[16'h0FA8] = 8'h00;
RAM[16'h0FA9] = 8'h00;
RAM[16'h0FAA] = 8'h00;
RAM[16'h0FAB] = 8'h00;
RAM[16'h0FAC] = 8'h00;
RAM[16'h0FAD] = 8'h00;
RAM[16'h0FAE] = 8'h00;
RAM[16'h0FAF] = 8'h00;
RAM[16'h0FB0] = 8'h00;
RAM[16'h0FB1] = 8'h00;
RAM[16'h0FB2] = 8'h00;
RAM[16'h0FB3] = 8'h00;
RAM[16'h0FB4] = 8'h00;
RAM[16'h0FB5] = 8'h00;
RAM[16'h0FB6] = 8'h00;
RAM[16'h0FB7] = 8'h00;
RAM[16'h0FB8] = 8'h00;
RAM[16'h0FB9] = 8'h00;
RAM[16'h0FBA] = 8'h00;
RAM[16'h0FBB] = 8'h00;
RAM[16'h0FBC] = 8'h00;
RAM[16'h0FBD] = 8'h00;
RAM[16'h0FBE] = 8'h00;
RAM[16'h0FBF] = 8'h00;
RAM[16'h0FC0] = 8'h00;
RAM[16'h0FC1] = 8'h00;
RAM[16'h0FC2] = 8'h00;
RAM[16'h0FC3] = 8'h00;
RAM[16'h0FC4] = 8'h00;
RAM[16'h0FC5] = 8'h00;
RAM[16'h0FC6] = 8'h00;
RAM[16'h0FC7] = 8'h00;
RAM[16'h0FC8] = 8'h00;
RAM[16'h0FC9] = 8'h00;
RAM[16'h0FCA] = 8'h00;
RAM[16'h0FCB] = 8'h00;
RAM[16'h0FCC] = 8'h00;
RAM[16'h0FCD] = 8'h00;
RAM[16'h0FCE] = 8'h00;
RAM[16'h0FCF] = 8'h00;
RAM[16'h0FD0] = 8'h00;
RAM[16'h0FD1] = 8'h00;
RAM[16'h0FD2] = 8'h00;
RAM[16'h0FD3] = 8'h00;
RAM[16'h0FD4] = 8'h00;
RAM[16'h0FD5] = 8'h00;
RAM[16'h0FD6] = 8'h00;
RAM[16'h0FD7] = 8'h00;
RAM[16'h0FD8] = 8'h00;
RAM[16'h0FD9] = 8'h00;
RAM[16'h0FDA] = 8'h00;
RAM[16'h0FDB] = 8'h00;
RAM[16'h0FDC] = 8'h00;
RAM[16'h0FDD] = 8'h00;
RAM[16'h0FDE] = 8'h00;
RAM[16'h0FDF] = 8'h00;
RAM[16'h0FE0] = 8'h00;
RAM[16'h0FE1] = 8'h00;
RAM[16'h0FE2] = 8'h00;
RAM[16'h0FE3] = 8'h00;
RAM[16'h0FE4] = 8'h00;
RAM[16'h0FE5] = 8'h00;
RAM[16'h0FE6] = 8'h00;
RAM[16'h0FE7] = 8'h00;
RAM[16'h0FE8] = 8'h00;
RAM[16'h0FE9] = 8'h00;
RAM[16'h0FEA] = 8'h00;
RAM[16'h0FEB] = 8'h00;
RAM[16'h0FEC] = 8'h00;
RAM[16'h0FED] = 8'h00;
RAM[16'h0FEE] = 8'h00;
RAM[16'h0FEF] = 8'h00;
RAM[16'h0FF0] = 8'h00;
RAM[16'h0FF1] = 8'h00;
RAM[16'h0FF2] = 8'h00;
RAM[16'h0FF3] = 8'h00;
RAM[16'h0FF4] = 8'h00;
RAM[16'h0FF5] = 8'h00;
RAM[16'h0FF6] = 8'h00;
RAM[16'h0FF7] = 8'h00;
RAM[16'h0FF8] = 8'h00;
RAM[16'h0FF9] = 8'h00;
RAM[16'h0FFA] = 8'h00;
RAM[16'h0FFB] = 8'h00;
RAM[16'h0FFC] = 8'h00;
RAM[16'h0FFD] = 8'h00;
RAM[16'h0FFE] = 8'h00;
RAM[16'h0FFF] = 8'h00;
RAM[16'h1000] = 8'h00;
RAM[16'h1001] = 8'h00;
RAM[16'h1002] = 8'h00;
RAM[16'h1003] = 8'h00;
RAM[16'h1004] = 8'h00;
RAM[16'h1005] = 8'h00;
RAM[16'h1006] = 8'h00;
RAM[16'h1007] = 8'h00;
RAM[16'h1008] = 8'h00;
RAM[16'h1009] = 8'h00;
RAM[16'h100A] = 8'h00;
RAM[16'h100B] = 8'h00;
RAM[16'h100C] = 8'h00;
RAM[16'h100D] = 8'h00;
RAM[16'h100E] = 8'h00;
RAM[16'h100F] = 8'h00;
RAM[16'h1010] = 8'h00;
RAM[16'h1011] = 8'h00;
RAM[16'h1012] = 8'h00;
RAM[16'h1013] = 8'h00;
RAM[16'h1014] = 8'h00;
RAM[16'h1015] = 8'h00;
RAM[16'h1016] = 8'h00;
RAM[16'h1017] = 8'h00;
RAM[16'h1018] = 8'h00;
RAM[16'h1019] = 8'h00;
RAM[16'h101A] = 8'h00;
RAM[16'h101B] = 8'h00;
RAM[16'h101C] = 8'h00;
RAM[16'h101D] = 8'h00;
RAM[16'h101E] = 8'h00;
RAM[16'h101F] = 8'h00;
RAM[16'h1020] = 8'h00;
RAM[16'h1021] = 8'h00;
RAM[16'h1022] = 8'h00;
RAM[16'h1023] = 8'h00;
RAM[16'h1024] = 8'h00;
RAM[16'h1025] = 8'h00;
RAM[16'h1026] = 8'h00;
RAM[16'h1027] = 8'h00;
RAM[16'h1028] = 8'h00;
RAM[16'h1029] = 8'h00;
RAM[16'h102A] = 8'h00;
RAM[16'h102B] = 8'h00;
RAM[16'h102C] = 8'h00;
RAM[16'h102D] = 8'h00;
RAM[16'h102E] = 8'h00;
RAM[16'h102F] = 8'h00;
RAM[16'h1030] = 8'h00;
RAM[16'h1031] = 8'h00;
RAM[16'h1032] = 8'h00;
RAM[16'h1033] = 8'h00;
RAM[16'h1034] = 8'h00;
RAM[16'h1035] = 8'h00;
RAM[16'h1036] = 8'h00;
RAM[16'h1037] = 8'h00;
RAM[16'h1038] = 8'h00;
RAM[16'h1039] = 8'h00;
RAM[16'h103A] = 8'h00;
RAM[16'h103B] = 8'h00;
RAM[16'h103C] = 8'h00;
RAM[16'h103D] = 8'h00;
RAM[16'h103E] = 8'h00;
RAM[16'h103F] = 8'h00;
RAM[16'h1040] = 8'h00;
RAM[16'h1041] = 8'h00;
RAM[16'h1042] = 8'h00;
RAM[16'h1043] = 8'h00;
RAM[16'h1044] = 8'h00;
RAM[16'h1045] = 8'h00;
RAM[16'h1046] = 8'h00;
RAM[16'h1047] = 8'h00;
RAM[16'h1048] = 8'h00;
RAM[16'h1049] = 8'h00;
RAM[16'h104A] = 8'h00;
RAM[16'h104B] = 8'h00;
RAM[16'h104C] = 8'h00;
RAM[16'h104D] = 8'h00;
RAM[16'h104E] = 8'h00;
RAM[16'h104F] = 8'h00;
RAM[16'h1050] = 8'h00;
RAM[16'h1051] = 8'h00;
RAM[16'h1052] = 8'h00;
RAM[16'h1053] = 8'h00;
RAM[16'h1054] = 8'h00;
RAM[16'h1055] = 8'h00;
RAM[16'h1056] = 8'h00;
RAM[16'h1057] = 8'h00;
RAM[16'h1058] = 8'h00;
RAM[16'h1059] = 8'h00;
RAM[16'h105A] = 8'h00;
RAM[16'h105B] = 8'h00;
RAM[16'h105C] = 8'h00;
RAM[16'h105D] = 8'h00;
RAM[16'h105E] = 8'h00;
RAM[16'h105F] = 8'h00;
RAM[16'h1060] = 8'h00;
RAM[16'h1061] = 8'h00;
RAM[16'h1062] = 8'h00;
RAM[16'h1063] = 8'h00;
RAM[16'h1064] = 8'h00;
RAM[16'h1065] = 8'h00;
RAM[16'h1066] = 8'h00;
RAM[16'h1067] = 8'h00;
RAM[16'h1068] = 8'h00;
RAM[16'h1069] = 8'h00;
RAM[16'h106A] = 8'h00;
RAM[16'h106B] = 8'h00;
RAM[16'h106C] = 8'h00;
RAM[16'h106D] = 8'h00;
RAM[16'h106E] = 8'h00;
RAM[16'h106F] = 8'h00;
RAM[16'h1070] = 8'h00;
RAM[16'h1071] = 8'h00;
RAM[16'h1072] = 8'h00;
RAM[16'h1073] = 8'h00;
RAM[16'h1074] = 8'h00;
RAM[16'h1075] = 8'h00;
RAM[16'h1076] = 8'h00;
RAM[16'h1077] = 8'h00;
RAM[16'h1078] = 8'h00;
RAM[16'h1079] = 8'h00;
RAM[16'h107A] = 8'h00;
RAM[16'h107B] = 8'h00;
RAM[16'h107C] = 8'h00;
RAM[16'h107D] = 8'h00;
RAM[16'h107E] = 8'h00;
RAM[16'h107F] = 8'h00;
RAM[16'h1080] = 8'h00;
RAM[16'h1081] = 8'h00;
RAM[16'h1082] = 8'h00;
RAM[16'h1083] = 8'h00;
RAM[16'h1084] = 8'h00;
RAM[16'h1085] = 8'h00;
RAM[16'h1086] = 8'h00;
RAM[16'h1087] = 8'h00;
RAM[16'h1088] = 8'h00;
RAM[16'h1089] = 8'h00;
RAM[16'h108A] = 8'h00;
RAM[16'h108B] = 8'h00;
RAM[16'h108C] = 8'h00;
RAM[16'h108D] = 8'h00;
RAM[16'h108E] = 8'h00;
RAM[16'h108F] = 8'h00;
RAM[16'h1090] = 8'h00;
RAM[16'h1091] = 8'h00;
RAM[16'h1092] = 8'h00;
RAM[16'h1093] = 8'h00;
RAM[16'h1094] = 8'h00;
RAM[16'h1095] = 8'h00;
RAM[16'h1096] = 8'h00;
RAM[16'h1097] = 8'h00;
RAM[16'h1098] = 8'h00;
RAM[16'h1099] = 8'h00;
RAM[16'h109A] = 8'h00;
RAM[16'h109B] = 8'h00;
RAM[16'h109C] = 8'h00;
RAM[16'h109D] = 8'h00;
RAM[16'h109E] = 8'h00;
RAM[16'h109F] = 8'h00;
RAM[16'h10A0] = 8'h00;
RAM[16'h10A1] = 8'h00;
RAM[16'h10A2] = 8'h00;
RAM[16'h10A3] = 8'h00;
RAM[16'h10A4] = 8'h00;
RAM[16'h10A5] = 8'h00;
RAM[16'h10A6] = 8'h00;
RAM[16'h10A7] = 8'h00;
RAM[16'h10A8] = 8'h00;
RAM[16'h10A9] = 8'h00;
RAM[16'h10AA] = 8'h00;
RAM[16'h10AB] = 8'h00;
RAM[16'h10AC] = 8'h00;
RAM[16'h10AD] = 8'h00;
RAM[16'h10AE] = 8'h00;
RAM[16'h10AF] = 8'h00;
RAM[16'h10B0] = 8'h00;
RAM[16'h10B1] = 8'h00;
RAM[16'h10B2] = 8'h00;
RAM[16'h10B3] = 8'h00;
RAM[16'h10B4] = 8'h00;
RAM[16'h10B5] = 8'h00;
RAM[16'h10B6] = 8'h00;
RAM[16'h10B7] = 8'h00;
RAM[16'h10B8] = 8'h00;
RAM[16'h10B9] = 8'h00;
RAM[16'h10BA] = 8'h00;
RAM[16'h10BB] = 8'h00;
RAM[16'h10BC] = 8'h00;
RAM[16'h10BD] = 8'h00;
RAM[16'h10BE] = 8'h00;
RAM[16'h10BF] = 8'h00;
RAM[16'h10C0] = 8'h00;
RAM[16'h10C1] = 8'h00;
RAM[16'h10C2] = 8'h00;
RAM[16'h10C3] = 8'h00;
RAM[16'h10C4] = 8'h00;
RAM[16'h10C5] = 8'h00;
RAM[16'h10C6] = 8'h00;
RAM[16'h10C7] = 8'h00;
RAM[16'h10C8] = 8'h00;
RAM[16'h10C9] = 8'h00;
RAM[16'h10CA] = 8'h00;
RAM[16'h10CB] = 8'h00;
RAM[16'h10CC] = 8'h00;
RAM[16'h10CD] = 8'h00;
RAM[16'h10CE] = 8'h00;
RAM[16'h10CF] = 8'h00;
RAM[16'h10D0] = 8'h00;
RAM[16'h10D1] = 8'h00;
RAM[16'h10D2] = 8'h00;
RAM[16'h10D3] = 8'h00;
RAM[16'h10D4] = 8'h00;
RAM[16'h10D5] = 8'h00;
RAM[16'h10D6] = 8'h00;
RAM[16'h10D7] = 8'h00;
RAM[16'h10D8] = 8'h00;
RAM[16'h10D9] = 8'h00;
RAM[16'h10DA] = 8'h00;
RAM[16'h10DB] = 8'h00;
RAM[16'h10DC] = 8'h00;
RAM[16'h10DD] = 8'h00;
RAM[16'h10DE] = 8'h00;
RAM[16'h10DF] = 8'h00;
RAM[16'h10E0] = 8'h00;
RAM[16'h10E1] = 8'h00;
RAM[16'h10E2] = 8'h00;
RAM[16'h10E3] = 8'h00;
RAM[16'h10E4] = 8'h00;
RAM[16'h10E5] = 8'h00;
RAM[16'h10E6] = 8'h00;
RAM[16'h10E7] = 8'h00;
RAM[16'h10E8] = 8'h00;
RAM[16'h10E9] = 8'h00;
RAM[16'h10EA] = 8'h00;
RAM[16'h10EB] = 8'h00;
RAM[16'h10EC] = 8'h00;
RAM[16'h10ED] = 8'h00;
RAM[16'h10EE] = 8'h00;
RAM[16'h10EF] = 8'h00;
RAM[16'h10F0] = 8'h00;
RAM[16'h10F1] = 8'h00;
RAM[16'h10F2] = 8'h00;
RAM[16'h10F3] = 8'h00;
RAM[16'h10F4] = 8'h00;
RAM[16'h10F5] = 8'h00;
RAM[16'h10F6] = 8'h00;
RAM[16'h10F7] = 8'h00;
RAM[16'h10F8] = 8'h00;
RAM[16'h10F9] = 8'h00;
RAM[16'h10FA] = 8'h00;
RAM[16'h10FB] = 8'h00;
RAM[16'h10FC] = 8'h00;
RAM[16'h10FD] = 8'h00;
RAM[16'h10FE] = 8'h00;
RAM[16'h10FF] = 8'h00;
RAM[16'h1100] = 8'h00;
RAM[16'h1101] = 8'h00;
RAM[16'h1102] = 8'h00;
RAM[16'h1103] = 8'h00;
RAM[16'h1104] = 8'h00;
RAM[16'h1105] = 8'h00;
RAM[16'h1106] = 8'h00;
RAM[16'h1107] = 8'h00;
RAM[16'h1108] = 8'h00;
RAM[16'h1109] = 8'h00;
RAM[16'h110A] = 8'h00;
RAM[16'h110B] = 8'h00;
RAM[16'h110C] = 8'h00;
RAM[16'h110D] = 8'h00;
RAM[16'h110E] = 8'h00;
RAM[16'h110F] = 8'h00;
RAM[16'h1110] = 8'h00;
RAM[16'h1111] = 8'h00;
RAM[16'h1112] = 8'h00;
RAM[16'h1113] = 8'h00;
RAM[16'h1114] = 8'h00;
RAM[16'h1115] = 8'h00;
RAM[16'h1116] = 8'h00;
RAM[16'h1117] = 8'h00;
RAM[16'h1118] = 8'h00;
RAM[16'h1119] = 8'h00;
RAM[16'h111A] = 8'h00;
RAM[16'h111B] = 8'h00;
RAM[16'h111C] = 8'h00;
RAM[16'h111D] = 8'h00;
RAM[16'h111E] = 8'h00;
RAM[16'h111F] = 8'h00;
RAM[16'h1120] = 8'h00;
RAM[16'h1121] = 8'h00;
RAM[16'h1122] = 8'h00;
RAM[16'h1123] = 8'h00;
RAM[16'h1124] = 8'h00;
RAM[16'h1125] = 8'h00;
RAM[16'h1126] = 8'h00;
RAM[16'h1127] = 8'h00;
RAM[16'h1128] = 8'h00;
RAM[16'h1129] = 8'h00;
RAM[16'h112A] = 8'h00;
RAM[16'h112B] = 8'h00;
RAM[16'h112C] = 8'h00;
RAM[16'h112D] = 8'h00;
RAM[16'h112E] = 8'h00;
RAM[16'h112F] = 8'h00;
RAM[16'h1130] = 8'h00;
RAM[16'h1131] = 8'h00;
RAM[16'h1132] = 8'h00;
RAM[16'h1133] = 8'h00;
RAM[16'h1134] = 8'h00;
RAM[16'h1135] = 8'h00;
RAM[16'h1136] = 8'h00;
RAM[16'h1137] = 8'h00;
RAM[16'h1138] = 8'h00;
RAM[16'h1139] = 8'h00;
RAM[16'h113A] = 8'h00;
RAM[16'h113B] = 8'h00;
RAM[16'h113C] = 8'h00;
RAM[16'h113D] = 8'h00;
RAM[16'h113E] = 8'h00;
RAM[16'h113F] = 8'h00;
RAM[16'h1140] = 8'h00;
RAM[16'h1141] = 8'h00;
RAM[16'h1142] = 8'h00;
RAM[16'h1143] = 8'h00;
RAM[16'h1144] = 8'h00;
RAM[16'h1145] = 8'h00;
RAM[16'h1146] = 8'h00;
RAM[16'h1147] = 8'h00;
RAM[16'h1148] = 8'h00;
RAM[16'h1149] = 8'h00;
RAM[16'h114A] = 8'h00;
RAM[16'h114B] = 8'h00;
RAM[16'h114C] = 8'h00;
RAM[16'h114D] = 8'h00;
RAM[16'h114E] = 8'h00;
RAM[16'h114F] = 8'h00;
RAM[16'h1150] = 8'h00;
RAM[16'h1151] = 8'h00;
RAM[16'h1152] = 8'h00;
RAM[16'h1153] = 8'h00;
RAM[16'h1154] = 8'h00;
RAM[16'h1155] = 8'h00;
RAM[16'h1156] = 8'h00;
RAM[16'h1157] = 8'h00;
RAM[16'h1158] = 8'h00;
RAM[16'h1159] = 8'h00;
RAM[16'h115A] = 8'h00;
RAM[16'h115B] = 8'h00;
RAM[16'h115C] = 8'h00;
RAM[16'h115D] = 8'h00;
RAM[16'h115E] = 8'h00;
RAM[16'h115F] = 8'h00;
RAM[16'h1160] = 8'h00;
RAM[16'h1161] = 8'h00;
RAM[16'h1162] = 8'h00;
RAM[16'h1163] = 8'h00;
RAM[16'h1164] = 8'h00;
RAM[16'h1165] = 8'h00;
RAM[16'h1166] = 8'h00;
RAM[16'h1167] = 8'h00;
RAM[16'h1168] = 8'h00;
RAM[16'h1169] = 8'h00;
RAM[16'h116A] = 8'h00;
RAM[16'h116B] = 8'h00;
RAM[16'h116C] = 8'h00;
RAM[16'h116D] = 8'h00;
RAM[16'h116E] = 8'h00;
RAM[16'h116F] = 8'h00;
RAM[16'h1170] = 8'h00;
RAM[16'h1171] = 8'h00;
RAM[16'h1172] = 8'h00;
RAM[16'h1173] = 8'h00;
RAM[16'h1174] = 8'h00;
RAM[16'h1175] = 8'h00;
RAM[16'h1176] = 8'h00;
RAM[16'h1177] = 8'h00;
RAM[16'h1178] = 8'h00;
RAM[16'h1179] = 8'h00;
RAM[16'h117A] = 8'h00;
RAM[16'h117B] = 8'h00;
RAM[16'h117C] = 8'h00;
RAM[16'h117D] = 8'h00;
RAM[16'h117E] = 8'h00;
RAM[16'h117F] = 8'h00;
RAM[16'h1180] = 8'h00;
RAM[16'h1181] = 8'h00;
RAM[16'h1182] = 8'h00;
RAM[16'h1183] = 8'h00;
RAM[16'h1184] = 8'h00;
RAM[16'h1185] = 8'h00;
RAM[16'h1186] = 8'h00;
RAM[16'h1187] = 8'h00;
RAM[16'h1188] = 8'h00;
RAM[16'h1189] = 8'h00;
RAM[16'h118A] = 8'h00;
RAM[16'h118B] = 8'h00;
RAM[16'h118C] = 8'h00;
RAM[16'h118D] = 8'h00;
RAM[16'h118E] = 8'h00;
RAM[16'h118F] = 8'h00;
RAM[16'h1190] = 8'h00;
RAM[16'h1191] = 8'h00;
RAM[16'h1192] = 8'h00;
RAM[16'h1193] = 8'h00;
RAM[16'h1194] = 8'h00;
RAM[16'h1195] = 8'h00;
RAM[16'h1196] = 8'h00;
RAM[16'h1197] = 8'h00;
RAM[16'h1198] = 8'h00;
RAM[16'h1199] = 8'h00;
RAM[16'h119A] = 8'h00;
RAM[16'h119B] = 8'h00;
RAM[16'h119C] = 8'h00;
RAM[16'h119D] = 8'h00;
RAM[16'h119E] = 8'h00;
RAM[16'h119F] = 8'h00;
RAM[16'h11A0] = 8'h00;
RAM[16'h11A1] = 8'h00;
RAM[16'h11A2] = 8'h00;
RAM[16'h11A3] = 8'h00;
RAM[16'h11A4] = 8'h00;
RAM[16'h11A5] = 8'h00;
RAM[16'h11A6] = 8'h00;
RAM[16'h11A7] = 8'h00;
RAM[16'h11A8] = 8'h00;
RAM[16'h11A9] = 8'h00;
RAM[16'h11AA] = 8'h00;
RAM[16'h11AB] = 8'h00;
RAM[16'h11AC] = 8'h00;
RAM[16'h11AD] = 8'h00;
RAM[16'h11AE] = 8'h00;
RAM[16'h11AF] = 8'h00;
RAM[16'h11B0] = 8'h00;
RAM[16'h11B1] = 8'h00;
RAM[16'h11B2] = 8'h00;
RAM[16'h11B3] = 8'h00;
RAM[16'h11B4] = 8'h00;
RAM[16'h11B5] = 8'h00;
RAM[16'h11B6] = 8'h00;
RAM[16'h11B7] = 8'h00;
RAM[16'h11B8] = 8'h00;
RAM[16'h11B9] = 8'h00;
RAM[16'h11BA] = 8'h00;
RAM[16'h11BB] = 8'h00;
RAM[16'h11BC] = 8'h00;
RAM[16'h11BD] = 8'h00;
RAM[16'h11BE] = 8'h00;
RAM[16'h11BF] = 8'h00;
RAM[16'h11C0] = 8'h00;
RAM[16'h11C1] = 8'h00;
RAM[16'h11C2] = 8'h00;
RAM[16'h11C3] = 8'h00;
RAM[16'h11C4] = 8'h00;
RAM[16'h11C5] = 8'h00;
RAM[16'h11C6] = 8'h00;
RAM[16'h11C7] = 8'h00;
RAM[16'h11C8] = 8'h00;
RAM[16'h11C9] = 8'h00;
RAM[16'h11CA] = 8'h00;
RAM[16'h11CB] = 8'h00;
RAM[16'h11CC] = 8'h00;
RAM[16'h11CD] = 8'h00;
RAM[16'h11CE] = 8'h00;
RAM[16'h11CF] = 8'h00;
RAM[16'h11D0] = 8'h00;
RAM[16'h11D1] = 8'h00;
RAM[16'h11D2] = 8'h00;
RAM[16'h11D3] = 8'h00;
RAM[16'h11D4] = 8'h00;
RAM[16'h11D5] = 8'h00;
RAM[16'h11D6] = 8'h00;
RAM[16'h11D7] = 8'h00;
RAM[16'h11D8] = 8'h00;
RAM[16'h11D9] = 8'h00;
RAM[16'h11DA] = 8'h00;
RAM[16'h11DB] = 8'h00;
RAM[16'h11DC] = 8'h00;
RAM[16'h11DD] = 8'h00;
RAM[16'h11DE] = 8'h00;
RAM[16'h11DF] = 8'h00;
RAM[16'h11E0] = 8'h00;
RAM[16'h11E1] = 8'h00;
RAM[16'h11E2] = 8'h00;
RAM[16'h11E3] = 8'h00;
RAM[16'h11E4] = 8'h00;
RAM[16'h11E5] = 8'h00;
RAM[16'h11E6] = 8'h00;
RAM[16'h11E7] = 8'h00;
RAM[16'h11E8] = 8'h00;
RAM[16'h11E9] = 8'h00;
RAM[16'h11EA] = 8'h00;
RAM[16'h11EB] = 8'h00;
RAM[16'h11EC] = 8'h00;
RAM[16'h11ED] = 8'h00;
RAM[16'h11EE] = 8'h00;
RAM[16'h11EF] = 8'h00;
RAM[16'h11F0] = 8'h00;
RAM[16'h11F1] = 8'h00;
RAM[16'h11F2] = 8'h00;
RAM[16'h11F3] = 8'h00;
RAM[16'h11F4] = 8'h00;
RAM[16'h11F5] = 8'h00;
RAM[16'h11F6] = 8'h00;
RAM[16'h11F7] = 8'h00;
RAM[16'h11F8] = 8'h00;
RAM[16'h11F9] = 8'h00;
RAM[16'h11FA] = 8'h00;
RAM[16'h11FB] = 8'h00;
RAM[16'h11FC] = 8'h00;
RAM[16'h11FD] = 8'h00;
RAM[16'h11FE] = 8'h00;
RAM[16'h11FF] = 8'h00;
RAM[16'h1200] = 8'h00;
RAM[16'h1201] = 8'h00;
RAM[16'h1202] = 8'h00;
RAM[16'h1203] = 8'h00;
RAM[16'h1204] = 8'h00;
RAM[16'h1205] = 8'h00;
RAM[16'h1206] = 8'h00;
RAM[16'h1207] = 8'h00;
RAM[16'h1208] = 8'h00;
RAM[16'h1209] = 8'h00;
RAM[16'h120A] = 8'h00;
RAM[16'h120B] = 8'h00;
RAM[16'h120C] = 8'h00;
RAM[16'h120D] = 8'h00;
RAM[16'h120E] = 8'h00;
RAM[16'h120F] = 8'h00;
RAM[16'h1210] = 8'h00;
RAM[16'h1211] = 8'h00;
RAM[16'h1212] = 8'h00;
RAM[16'h1213] = 8'h00;
RAM[16'h1214] = 8'h00;
RAM[16'h1215] = 8'h00;
RAM[16'h1216] = 8'h00;
RAM[16'h1217] = 8'h00;
RAM[16'h1218] = 8'h00;
RAM[16'h1219] = 8'h00;
RAM[16'h121A] = 8'h00;
RAM[16'h121B] = 8'h00;
RAM[16'h121C] = 8'h00;
RAM[16'h121D] = 8'h00;
RAM[16'h121E] = 8'h00;
RAM[16'h121F] = 8'h00;
RAM[16'h1220] = 8'h00;
RAM[16'h1221] = 8'h00;
RAM[16'h1222] = 8'h00;
RAM[16'h1223] = 8'h00;
RAM[16'h1224] = 8'h00;
RAM[16'h1225] = 8'h00;
RAM[16'h1226] = 8'h00;
RAM[16'h1227] = 8'h00;
RAM[16'h1228] = 8'h00;
RAM[16'h1229] = 8'h00;
RAM[16'h122A] = 8'h00;
RAM[16'h122B] = 8'h00;
RAM[16'h122C] = 8'h00;
RAM[16'h122D] = 8'h00;
RAM[16'h122E] = 8'h00;
RAM[16'h122F] = 8'h00;
RAM[16'h1230] = 8'h00;
RAM[16'h1231] = 8'h00;
RAM[16'h1232] = 8'h00;
RAM[16'h1233] = 8'h00;
RAM[16'h1234] = 8'h00;
RAM[16'h1235] = 8'h00;
RAM[16'h1236] = 8'h00;
RAM[16'h1237] = 8'h00;
RAM[16'h1238] = 8'h00;
RAM[16'h1239] = 8'h00;
RAM[16'h123A] = 8'h00;
RAM[16'h123B] = 8'h00;
RAM[16'h123C] = 8'h00;
RAM[16'h123D] = 8'h00;
RAM[16'h123E] = 8'h00;
RAM[16'h123F] = 8'h00;
RAM[16'h1240] = 8'h00;
RAM[16'h1241] = 8'h00;
RAM[16'h1242] = 8'h00;
RAM[16'h1243] = 8'h00;
RAM[16'h1244] = 8'h00;
RAM[16'h1245] = 8'h00;
RAM[16'h1246] = 8'h00;
RAM[16'h1247] = 8'h00;
RAM[16'h1248] = 8'h00;
RAM[16'h1249] = 8'h00;
RAM[16'h124A] = 8'h00;
RAM[16'h124B] = 8'h00;
RAM[16'h124C] = 8'h00;
RAM[16'h124D] = 8'h00;
RAM[16'h124E] = 8'h00;
RAM[16'h124F] = 8'h00;
RAM[16'h1250] = 8'h00;
RAM[16'h1251] = 8'h00;
RAM[16'h1252] = 8'h00;
RAM[16'h1253] = 8'h00;
RAM[16'h1254] = 8'h00;
RAM[16'h1255] = 8'h00;
RAM[16'h1256] = 8'h00;
RAM[16'h1257] = 8'h00;
RAM[16'h1258] = 8'h00;
RAM[16'h1259] = 8'h00;
RAM[16'h125A] = 8'h00;
RAM[16'h125B] = 8'h00;
RAM[16'h125C] = 8'h00;
RAM[16'h125D] = 8'h00;
RAM[16'h125E] = 8'h00;
RAM[16'h125F] = 8'h00;
RAM[16'h1260] = 8'h00;
RAM[16'h1261] = 8'h00;
RAM[16'h1262] = 8'h00;
RAM[16'h1263] = 8'h00;
RAM[16'h1264] = 8'h00;
RAM[16'h1265] = 8'h00;
RAM[16'h1266] = 8'h00;
RAM[16'h1267] = 8'h00;
RAM[16'h1268] = 8'h00;
RAM[16'h1269] = 8'h00;
RAM[16'h126A] = 8'h00;
RAM[16'h126B] = 8'h00;
RAM[16'h126C] = 8'h00;
RAM[16'h126D] = 8'h00;
RAM[16'h126E] = 8'h00;
RAM[16'h126F] = 8'h00;
RAM[16'h1270] = 8'h00;
RAM[16'h1271] = 8'h00;
RAM[16'h1272] = 8'h00;
RAM[16'h1273] = 8'h00;
RAM[16'h1274] = 8'h00;
RAM[16'h1275] = 8'h00;
RAM[16'h1276] = 8'h00;
RAM[16'h1277] = 8'h00;
RAM[16'h1278] = 8'h00;
RAM[16'h1279] = 8'h00;
RAM[16'h127A] = 8'h00;
RAM[16'h127B] = 8'h00;
RAM[16'h127C] = 8'h00;
RAM[16'h127D] = 8'h00;
RAM[16'h127E] = 8'h00;
RAM[16'h127F] = 8'h00;
RAM[16'h1280] = 8'h00;
RAM[16'h1281] = 8'h00;
RAM[16'h1282] = 8'h00;
RAM[16'h1283] = 8'h00;
RAM[16'h1284] = 8'h00;
RAM[16'h1285] = 8'h00;
RAM[16'h1286] = 8'h00;
RAM[16'h1287] = 8'h00;
RAM[16'h1288] = 8'h00;
RAM[16'h1289] = 8'h00;
RAM[16'h128A] = 8'h00;
RAM[16'h128B] = 8'h00;
RAM[16'h128C] = 8'h00;
RAM[16'h128D] = 8'h00;
RAM[16'h128E] = 8'h00;
RAM[16'h128F] = 8'h00;
RAM[16'h1290] = 8'h00;
RAM[16'h1291] = 8'h00;
RAM[16'h1292] = 8'h00;
RAM[16'h1293] = 8'h00;
RAM[16'h1294] = 8'h00;
RAM[16'h1295] = 8'h00;
RAM[16'h1296] = 8'h00;
RAM[16'h1297] = 8'h00;
RAM[16'h1298] = 8'h00;
RAM[16'h1299] = 8'h00;
RAM[16'h129A] = 8'h00;
RAM[16'h129B] = 8'h00;
RAM[16'h129C] = 8'h00;
RAM[16'h129D] = 8'h00;
RAM[16'h129E] = 8'h00;
RAM[16'h129F] = 8'h00;
RAM[16'h12A0] = 8'h00;
RAM[16'h12A1] = 8'h00;
RAM[16'h12A2] = 8'h00;
RAM[16'h12A3] = 8'h00;
RAM[16'h12A4] = 8'h00;
RAM[16'h12A5] = 8'h00;
RAM[16'h12A6] = 8'h00;
RAM[16'h12A7] = 8'h00;
RAM[16'h12A8] = 8'h00;
RAM[16'h12A9] = 8'h00;
RAM[16'h12AA] = 8'h00;
RAM[16'h12AB] = 8'h00;
RAM[16'h12AC] = 8'h00;
RAM[16'h12AD] = 8'h00;
RAM[16'h12AE] = 8'h00;
RAM[16'h12AF] = 8'h00;
RAM[16'h12B0] = 8'h00;
RAM[16'h12B1] = 8'h00;
RAM[16'h12B2] = 8'h00;
RAM[16'h12B3] = 8'h00;
RAM[16'h12B4] = 8'h00;
RAM[16'h12B5] = 8'h00;
RAM[16'h12B6] = 8'h00;
RAM[16'h12B7] = 8'h00;
RAM[16'h12B8] = 8'h00;
RAM[16'h12B9] = 8'h00;
RAM[16'h12BA] = 8'h00;
RAM[16'h12BB] = 8'h00;
RAM[16'h12BC] = 8'h00;
RAM[16'h12BD] = 8'h00;
RAM[16'h12BE] = 8'h00;
RAM[16'h12BF] = 8'h00;
RAM[16'h12C0] = 8'h00;
RAM[16'h12C1] = 8'h00;
RAM[16'h12C2] = 8'h00;
RAM[16'h12C3] = 8'h00;
RAM[16'h12C4] = 8'h00;
RAM[16'h12C5] = 8'h00;
RAM[16'h12C6] = 8'h00;
RAM[16'h12C7] = 8'h00;
RAM[16'h12C8] = 8'h00;
RAM[16'h12C9] = 8'h00;
RAM[16'h12CA] = 8'h00;
RAM[16'h12CB] = 8'h00;
RAM[16'h12CC] = 8'h00;
RAM[16'h12CD] = 8'h00;
RAM[16'h12CE] = 8'h00;
RAM[16'h12CF] = 8'h00;
RAM[16'h12D0] = 8'h00;
RAM[16'h12D1] = 8'h00;
RAM[16'h12D2] = 8'h00;
RAM[16'h12D3] = 8'h00;
RAM[16'h12D4] = 8'h00;
RAM[16'h12D5] = 8'h00;
RAM[16'h12D6] = 8'h00;
RAM[16'h12D7] = 8'h00;
RAM[16'h12D8] = 8'h00;
RAM[16'h12D9] = 8'h00;
RAM[16'h12DA] = 8'h00;
RAM[16'h12DB] = 8'h00;
RAM[16'h12DC] = 8'h00;
RAM[16'h12DD] = 8'h00;
RAM[16'h12DE] = 8'h00;
RAM[16'h12DF] = 8'h00;
RAM[16'h12E0] = 8'h00;
RAM[16'h12E1] = 8'h00;
RAM[16'h12E2] = 8'h00;
RAM[16'h12E3] = 8'h00;
RAM[16'h12E4] = 8'h00;
RAM[16'h12E5] = 8'h00;
RAM[16'h12E6] = 8'h00;
RAM[16'h12E7] = 8'h00;
RAM[16'h12E8] = 8'h00;
RAM[16'h12E9] = 8'h00;
RAM[16'h12EA] = 8'h00;
RAM[16'h12EB] = 8'h00;
RAM[16'h12EC] = 8'h00;
RAM[16'h12ED] = 8'h00;
RAM[16'h12EE] = 8'h00;
RAM[16'h12EF] = 8'h00;
RAM[16'h12F0] = 8'h00;
RAM[16'h12F1] = 8'h00;
RAM[16'h12F2] = 8'h00;
RAM[16'h12F3] = 8'h00;
RAM[16'h12F4] = 8'h00;
RAM[16'h12F5] = 8'h00;
RAM[16'h12F6] = 8'h00;
RAM[16'h12F7] = 8'h00;
RAM[16'h12F8] = 8'h00;
RAM[16'h12F9] = 8'h00;
RAM[16'h12FA] = 8'h00;
RAM[16'h12FB] = 8'h00;
RAM[16'h12FC] = 8'h00;
RAM[16'h12FD] = 8'h00;
RAM[16'h12FE] = 8'h00;
RAM[16'h12FF] = 8'h00;
RAM[16'h1300] = 8'h00;
RAM[16'h1301] = 8'h00;
RAM[16'h1302] = 8'h00;
RAM[16'h1303] = 8'h00;
RAM[16'h1304] = 8'h00;
RAM[16'h1305] = 8'h00;
RAM[16'h1306] = 8'h00;
RAM[16'h1307] = 8'h00;
RAM[16'h1308] = 8'h00;
RAM[16'h1309] = 8'h00;
RAM[16'h130A] = 8'h00;
RAM[16'h130B] = 8'h00;
RAM[16'h130C] = 8'h00;
RAM[16'h130D] = 8'h00;
RAM[16'h130E] = 8'h00;
RAM[16'h130F] = 8'h00;
RAM[16'h1310] = 8'h00;
RAM[16'h1311] = 8'h00;
RAM[16'h1312] = 8'h00;
RAM[16'h1313] = 8'h00;
RAM[16'h1314] = 8'h00;
RAM[16'h1315] = 8'h00;
RAM[16'h1316] = 8'h00;
RAM[16'h1317] = 8'h00;
RAM[16'h1318] = 8'h00;
RAM[16'h1319] = 8'h00;
RAM[16'h131A] = 8'h00;
RAM[16'h131B] = 8'h00;
RAM[16'h131C] = 8'h00;
RAM[16'h131D] = 8'h00;
RAM[16'h131E] = 8'h00;
RAM[16'h131F] = 8'h00;
RAM[16'h1320] = 8'h00;
RAM[16'h1321] = 8'h00;
RAM[16'h1322] = 8'h00;
RAM[16'h1323] = 8'h00;
RAM[16'h1324] = 8'h00;
RAM[16'h1325] = 8'h00;
RAM[16'h1326] = 8'h00;
RAM[16'h1327] = 8'h00;
RAM[16'h1328] = 8'h00;
RAM[16'h1329] = 8'h00;
RAM[16'h132A] = 8'h00;
RAM[16'h132B] = 8'h00;
RAM[16'h132C] = 8'h00;
RAM[16'h132D] = 8'h00;
RAM[16'h132E] = 8'h00;
RAM[16'h132F] = 8'h00;
RAM[16'h1330] = 8'h00;
RAM[16'h1331] = 8'h00;
RAM[16'h1332] = 8'h00;
RAM[16'h1333] = 8'h00;
RAM[16'h1334] = 8'h00;
RAM[16'h1335] = 8'h00;
RAM[16'h1336] = 8'h00;
RAM[16'h1337] = 8'h00;
RAM[16'h1338] = 8'h00;
RAM[16'h1339] = 8'h00;
RAM[16'h133A] = 8'h00;
RAM[16'h133B] = 8'h00;
RAM[16'h133C] = 8'h00;
RAM[16'h133D] = 8'h00;
RAM[16'h133E] = 8'h00;
RAM[16'h133F] = 8'h00;
RAM[16'h1340] = 8'h00;
RAM[16'h1341] = 8'h00;
RAM[16'h1342] = 8'h00;
RAM[16'h1343] = 8'h00;
RAM[16'h1344] = 8'h00;
RAM[16'h1345] = 8'h00;
RAM[16'h1346] = 8'h00;
RAM[16'h1347] = 8'h00;
RAM[16'h1348] = 8'h00;
RAM[16'h1349] = 8'h00;
RAM[16'h134A] = 8'h00;
RAM[16'h134B] = 8'h00;
RAM[16'h134C] = 8'h00;
RAM[16'h134D] = 8'h00;
RAM[16'h134E] = 8'h00;
RAM[16'h134F] = 8'h00;
RAM[16'h1350] = 8'h00;
RAM[16'h1351] = 8'h00;
RAM[16'h1352] = 8'h00;
RAM[16'h1353] = 8'h00;
RAM[16'h1354] = 8'h00;
RAM[16'h1355] = 8'h00;
RAM[16'h1356] = 8'h00;
RAM[16'h1357] = 8'h00;
RAM[16'h1358] = 8'h00;
RAM[16'h1359] = 8'h00;
RAM[16'h135A] = 8'h00;
RAM[16'h135B] = 8'h00;
RAM[16'h135C] = 8'h00;
RAM[16'h135D] = 8'h00;
RAM[16'h135E] = 8'h00;
RAM[16'h135F] = 8'h00;
RAM[16'h1360] = 8'h00;
RAM[16'h1361] = 8'h00;
RAM[16'h1362] = 8'h00;
RAM[16'h1363] = 8'h00;
RAM[16'h1364] = 8'h00;
RAM[16'h1365] = 8'h00;
RAM[16'h1366] = 8'h00;
RAM[16'h1367] = 8'h00;
RAM[16'h1368] = 8'h00;
RAM[16'h1369] = 8'h00;
RAM[16'h136A] = 8'h00;
RAM[16'h136B] = 8'h00;
RAM[16'h136C] = 8'h00;
RAM[16'h136D] = 8'h00;
RAM[16'h136E] = 8'h00;
RAM[16'h136F] = 8'h00;
RAM[16'h1370] = 8'h00;
RAM[16'h1371] = 8'h00;
RAM[16'h1372] = 8'h00;
RAM[16'h1373] = 8'h00;
RAM[16'h1374] = 8'h00;
RAM[16'h1375] = 8'h00;
RAM[16'h1376] = 8'h00;
RAM[16'h1377] = 8'h00;
RAM[16'h1378] = 8'h00;
RAM[16'h1379] = 8'h00;
RAM[16'h137A] = 8'h00;
RAM[16'h137B] = 8'h00;
RAM[16'h137C] = 8'h00;
RAM[16'h137D] = 8'h00;
RAM[16'h137E] = 8'h00;
RAM[16'h137F] = 8'h00;
RAM[16'h1380] = 8'h00;
RAM[16'h1381] = 8'h00;
RAM[16'h1382] = 8'h00;
RAM[16'h1383] = 8'h00;
RAM[16'h1384] = 8'h00;
RAM[16'h1385] = 8'h00;
RAM[16'h1386] = 8'h00;
RAM[16'h1387] = 8'h00;
RAM[16'h1388] = 8'h00;
RAM[16'h1389] = 8'h00;
RAM[16'h138A] = 8'h00;
RAM[16'h138B] = 8'h00;
RAM[16'h138C] = 8'h00;
RAM[16'h138D] = 8'h00;
RAM[16'h138E] = 8'h00;
RAM[16'h138F] = 8'h00;
RAM[16'h1390] = 8'h00;
RAM[16'h1391] = 8'h00;
RAM[16'h1392] = 8'h00;
RAM[16'h1393] = 8'h00;
RAM[16'h1394] = 8'h00;
RAM[16'h1395] = 8'h00;
RAM[16'h1396] = 8'h00;
RAM[16'h1397] = 8'h00;
RAM[16'h1398] = 8'h00;
RAM[16'h1399] = 8'h00;
RAM[16'h139A] = 8'h00;
RAM[16'h139B] = 8'h00;
RAM[16'h139C] = 8'h00;
RAM[16'h139D] = 8'h00;
RAM[16'h139E] = 8'h00;
RAM[16'h139F] = 8'h00;
RAM[16'h13A0] = 8'h00;
RAM[16'h13A1] = 8'h00;
RAM[16'h13A2] = 8'h00;
RAM[16'h13A3] = 8'h00;
RAM[16'h13A4] = 8'h00;
RAM[16'h13A5] = 8'h00;
RAM[16'h13A6] = 8'h00;
RAM[16'h13A7] = 8'h00;
RAM[16'h13A8] = 8'h00;
RAM[16'h13A9] = 8'h00;
RAM[16'h13AA] = 8'h00;
RAM[16'h13AB] = 8'h00;
RAM[16'h13AC] = 8'h00;
RAM[16'h13AD] = 8'h00;
RAM[16'h13AE] = 8'h00;
RAM[16'h13AF] = 8'h00;
RAM[16'h13B0] = 8'h00;
RAM[16'h13B1] = 8'h00;
RAM[16'h13B2] = 8'h00;
RAM[16'h13B3] = 8'h00;
RAM[16'h13B4] = 8'h00;
RAM[16'h13B5] = 8'h00;
RAM[16'h13B6] = 8'h00;
RAM[16'h13B7] = 8'h00;
RAM[16'h13B8] = 8'h00;
RAM[16'h13B9] = 8'h00;
RAM[16'h13BA] = 8'h00;
RAM[16'h13BB] = 8'h00;
RAM[16'h13BC] = 8'h00;
RAM[16'h13BD] = 8'h00;
RAM[16'h13BE] = 8'h00;
RAM[16'h13BF] = 8'h00;
RAM[16'h13C0] = 8'h00;
RAM[16'h13C1] = 8'h00;
RAM[16'h13C2] = 8'h00;
RAM[16'h13C3] = 8'h00;
RAM[16'h13C4] = 8'h00;
RAM[16'h13C5] = 8'h00;
RAM[16'h13C6] = 8'h00;
RAM[16'h13C7] = 8'h00;
RAM[16'h13C8] = 8'h00;
RAM[16'h13C9] = 8'h00;
RAM[16'h13CA] = 8'h00;
RAM[16'h13CB] = 8'h00;
RAM[16'h13CC] = 8'h00;
RAM[16'h13CD] = 8'h00;
RAM[16'h13CE] = 8'h00;
RAM[16'h13CF] = 8'h00;
RAM[16'h13D0] = 8'h00;
RAM[16'h13D1] = 8'h00;
RAM[16'h13D2] = 8'h00;
RAM[16'h13D3] = 8'h00;
RAM[16'h13D4] = 8'h00;
RAM[16'h13D5] = 8'h00;
RAM[16'h13D6] = 8'h00;
RAM[16'h13D7] = 8'h00;
RAM[16'h13D8] = 8'h00;
RAM[16'h13D9] = 8'h00;
RAM[16'h13DA] = 8'h00;
RAM[16'h13DB] = 8'h00;
RAM[16'h13DC] = 8'h00;
RAM[16'h13DD] = 8'h00;
RAM[16'h13DE] = 8'h00;
RAM[16'h13DF] = 8'h00;
RAM[16'h13E0] = 8'h00;
RAM[16'h13E1] = 8'h00;
RAM[16'h13E2] = 8'h00;
RAM[16'h13E3] = 8'h00;
RAM[16'h13E4] = 8'h00;
RAM[16'h13E5] = 8'h00;
RAM[16'h13E6] = 8'h00;
RAM[16'h13E7] = 8'h00;
RAM[16'h13E8] = 8'h00;
RAM[16'h13E9] = 8'h00;
RAM[16'h13EA] = 8'h00;
RAM[16'h13EB] = 8'h00;
RAM[16'h13EC] = 8'h00;
RAM[16'h13ED] = 8'h00;
RAM[16'h13EE] = 8'h00;
RAM[16'h13EF] = 8'h00;
RAM[16'h13F0] = 8'h00;
RAM[16'h13F1] = 8'h00;
RAM[16'h13F2] = 8'h00;
RAM[16'h13F3] = 8'h00;
RAM[16'h13F4] = 8'h00;
RAM[16'h13F5] = 8'h00;
RAM[16'h13F6] = 8'h00;
RAM[16'h13F7] = 8'h00;
RAM[16'h13F8] = 8'h00;
RAM[16'h13F9] = 8'h00;
RAM[16'h13FA] = 8'h00;
RAM[16'h13FB] = 8'h00;
RAM[16'h13FC] = 8'h00;
RAM[16'h13FD] = 8'h00;
RAM[16'h13FE] = 8'h00;
RAM[16'h13FF] = 8'h00;
RAM[16'h1400] = 8'h00;
RAM[16'h1401] = 8'h00;
RAM[16'h1402] = 8'h00;
RAM[16'h1403] = 8'h00;
RAM[16'h1404] = 8'h00;
RAM[16'h1405] = 8'h00;
RAM[16'h1406] = 8'h00;
RAM[16'h1407] = 8'h00;
RAM[16'h1408] = 8'h00;
RAM[16'h1409] = 8'h00;
RAM[16'h140A] = 8'h00;
RAM[16'h140B] = 8'h00;
RAM[16'h140C] = 8'h00;
RAM[16'h140D] = 8'h00;
RAM[16'h140E] = 8'h00;
RAM[16'h140F] = 8'h00;
RAM[16'h1410] = 8'h00;
RAM[16'h1411] = 8'h00;
RAM[16'h1412] = 8'h00;
RAM[16'h1413] = 8'h00;
RAM[16'h1414] = 8'h00;
RAM[16'h1415] = 8'h00;
RAM[16'h1416] = 8'h00;
RAM[16'h1417] = 8'h00;
RAM[16'h1418] = 8'h00;
RAM[16'h1419] = 8'h00;
RAM[16'h141A] = 8'h00;
RAM[16'h141B] = 8'h00;
RAM[16'h141C] = 8'h00;
RAM[16'h141D] = 8'h00;
RAM[16'h141E] = 8'h00;
RAM[16'h141F] = 8'h00;
RAM[16'h1420] = 8'h00;
RAM[16'h1421] = 8'h00;
RAM[16'h1422] = 8'h00;
RAM[16'h1423] = 8'h00;
RAM[16'h1424] = 8'h00;
RAM[16'h1425] = 8'h00;
RAM[16'h1426] = 8'h00;
RAM[16'h1427] = 8'h00;
RAM[16'h1428] = 8'h00;
RAM[16'h1429] = 8'h00;
RAM[16'h142A] = 8'h00;
RAM[16'h142B] = 8'h00;
RAM[16'h142C] = 8'h00;
RAM[16'h142D] = 8'h00;
RAM[16'h142E] = 8'h00;
RAM[16'h142F] = 8'h00;
RAM[16'h1430] = 8'h00;
RAM[16'h1431] = 8'h00;
RAM[16'h1432] = 8'h00;
RAM[16'h1433] = 8'h00;
RAM[16'h1434] = 8'h00;
RAM[16'h1435] = 8'h00;
RAM[16'h1436] = 8'h00;
RAM[16'h1437] = 8'h00;
RAM[16'h1438] = 8'h00;
RAM[16'h1439] = 8'h00;
RAM[16'h143A] = 8'h00;
RAM[16'h143B] = 8'h00;
RAM[16'h143C] = 8'h00;
RAM[16'h143D] = 8'h00;
RAM[16'h143E] = 8'h00;
RAM[16'h143F] = 8'h00;
RAM[16'h1440] = 8'h00;
RAM[16'h1441] = 8'h00;
RAM[16'h1442] = 8'h00;
RAM[16'h1443] = 8'h00;
RAM[16'h1444] = 8'h00;
RAM[16'h1445] = 8'h00;
RAM[16'h1446] = 8'h00;
RAM[16'h1447] = 8'h00;
RAM[16'h1448] = 8'h00;
RAM[16'h1449] = 8'h00;
RAM[16'h144A] = 8'h00;
RAM[16'h144B] = 8'h00;
RAM[16'h144C] = 8'h00;
RAM[16'h144D] = 8'h00;
RAM[16'h144E] = 8'h00;
RAM[16'h144F] = 8'h00;
RAM[16'h1450] = 8'h00;
RAM[16'h1451] = 8'h00;
RAM[16'h1452] = 8'h00;
RAM[16'h1453] = 8'h00;
RAM[16'h1454] = 8'h00;
RAM[16'h1455] = 8'h00;
RAM[16'h1456] = 8'h00;
RAM[16'h1457] = 8'h00;
RAM[16'h1458] = 8'h00;
RAM[16'h1459] = 8'h00;
RAM[16'h145A] = 8'h00;
RAM[16'h145B] = 8'h00;
RAM[16'h145C] = 8'h00;
RAM[16'h145D] = 8'h00;
RAM[16'h145E] = 8'h00;
RAM[16'h145F] = 8'h00;
RAM[16'h1460] = 8'h00;
RAM[16'h1461] = 8'h00;
RAM[16'h1462] = 8'h00;
RAM[16'h1463] = 8'h00;
RAM[16'h1464] = 8'h00;
RAM[16'h1465] = 8'h00;
RAM[16'h1466] = 8'h00;
RAM[16'h1467] = 8'h00;
RAM[16'h1468] = 8'h00;
RAM[16'h1469] = 8'h00;
RAM[16'h146A] = 8'h00;
RAM[16'h146B] = 8'h00;
RAM[16'h146C] = 8'h00;
RAM[16'h146D] = 8'h00;
RAM[16'h146E] = 8'h00;
RAM[16'h146F] = 8'h00;
RAM[16'h1470] = 8'h00;
RAM[16'h1471] = 8'h00;
RAM[16'h1472] = 8'h00;
RAM[16'h1473] = 8'h00;
RAM[16'h1474] = 8'h00;
RAM[16'h1475] = 8'h00;
RAM[16'h1476] = 8'h00;
RAM[16'h1477] = 8'h00;
RAM[16'h1478] = 8'h00;
RAM[16'h1479] = 8'h00;
RAM[16'h147A] = 8'h00;
RAM[16'h147B] = 8'h00;
RAM[16'h147C] = 8'h00;
RAM[16'h147D] = 8'h00;
RAM[16'h147E] = 8'h00;
RAM[16'h147F] = 8'h00;
RAM[16'h1480] = 8'h00;
RAM[16'h1481] = 8'h00;
RAM[16'h1482] = 8'h00;
RAM[16'h1483] = 8'h00;
RAM[16'h1484] = 8'h00;
RAM[16'h1485] = 8'h00;
RAM[16'h1486] = 8'h00;
RAM[16'h1487] = 8'h00;
RAM[16'h1488] = 8'h00;
RAM[16'h1489] = 8'h00;
RAM[16'h148A] = 8'h00;
RAM[16'h148B] = 8'h00;
RAM[16'h148C] = 8'h00;
RAM[16'h148D] = 8'h00;
RAM[16'h148E] = 8'h00;
RAM[16'h148F] = 8'h00;
RAM[16'h1490] = 8'h00;
RAM[16'h1491] = 8'h00;
RAM[16'h1492] = 8'h00;
RAM[16'h1493] = 8'h00;
RAM[16'h1494] = 8'h00;
RAM[16'h1495] = 8'h00;
RAM[16'h1496] = 8'h00;
RAM[16'h1497] = 8'h00;
RAM[16'h1498] = 8'h00;
RAM[16'h1499] = 8'h00;
RAM[16'h149A] = 8'h00;
RAM[16'h149B] = 8'h00;
RAM[16'h149C] = 8'h00;
RAM[16'h149D] = 8'h00;
RAM[16'h149E] = 8'h00;
RAM[16'h149F] = 8'h00;
RAM[16'h14A0] = 8'h00;
RAM[16'h14A1] = 8'h00;
RAM[16'h14A2] = 8'h00;
RAM[16'h14A3] = 8'h00;
RAM[16'h14A4] = 8'h00;
RAM[16'h14A5] = 8'h00;
RAM[16'h14A6] = 8'h00;
RAM[16'h14A7] = 8'h00;
RAM[16'h14A8] = 8'h00;
RAM[16'h14A9] = 8'h00;
RAM[16'h14AA] = 8'h00;
RAM[16'h14AB] = 8'h00;
RAM[16'h14AC] = 8'h00;
RAM[16'h14AD] = 8'h00;
RAM[16'h14AE] = 8'h00;
RAM[16'h14AF] = 8'h00;
RAM[16'h14B0] = 8'h00;
RAM[16'h14B1] = 8'h00;
RAM[16'h14B2] = 8'h00;
RAM[16'h14B3] = 8'h00;
RAM[16'h14B4] = 8'h00;
RAM[16'h14B5] = 8'h00;
RAM[16'h14B6] = 8'h00;
RAM[16'h14B7] = 8'h00;
RAM[16'h14B8] = 8'h00;
RAM[16'h14B9] = 8'h00;
RAM[16'h14BA] = 8'h00;
RAM[16'h14BB] = 8'h00;
RAM[16'h14BC] = 8'h00;
RAM[16'h14BD] = 8'h00;
RAM[16'h14BE] = 8'h00;
RAM[16'h14BF] = 8'h00;
RAM[16'h14C0] = 8'h00;
RAM[16'h14C1] = 8'h00;
RAM[16'h14C2] = 8'h00;
RAM[16'h14C3] = 8'h00;
RAM[16'h14C4] = 8'h00;
RAM[16'h14C5] = 8'h00;
RAM[16'h14C6] = 8'h00;
RAM[16'h14C7] = 8'h00;
RAM[16'h14C8] = 8'h00;
RAM[16'h14C9] = 8'h00;
RAM[16'h14CA] = 8'h00;
RAM[16'h14CB] = 8'h00;
RAM[16'h14CC] = 8'h00;
RAM[16'h14CD] = 8'h00;
RAM[16'h14CE] = 8'h00;
RAM[16'h14CF] = 8'h00;
RAM[16'h14D0] = 8'h00;
RAM[16'h14D1] = 8'h00;
RAM[16'h14D2] = 8'h00;
RAM[16'h14D3] = 8'h00;
RAM[16'h14D4] = 8'h00;
RAM[16'h14D5] = 8'h00;
RAM[16'h14D6] = 8'h00;
RAM[16'h14D7] = 8'h00;
RAM[16'h14D8] = 8'h00;
RAM[16'h14D9] = 8'h00;
RAM[16'h14DA] = 8'h00;
RAM[16'h14DB] = 8'h00;
RAM[16'h14DC] = 8'h00;
RAM[16'h14DD] = 8'h00;
RAM[16'h14DE] = 8'h00;
RAM[16'h14DF] = 8'h00;
RAM[16'h14E0] = 8'h00;
RAM[16'h14E1] = 8'h00;
RAM[16'h14E2] = 8'h00;
RAM[16'h14E3] = 8'h00;
RAM[16'h14E4] = 8'h00;
RAM[16'h14E5] = 8'h00;
RAM[16'h14E6] = 8'h00;
RAM[16'h14E7] = 8'h00;
RAM[16'h14E8] = 8'h00;
RAM[16'h14E9] = 8'h00;
RAM[16'h14EA] = 8'h00;
RAM[16'h14EB] = 8'h00;
RAM[16'h14EC] = 8'h00;
RAM[16'h14ED] = 8'h00;
RAM[16'h14EE] = 8'h00;
RAM[16'h14EF] = 8'h00;
RAM[16'h14F0] = 8'h00;
RAM[16'h14F1] = 8'h00;
RAM[16'h14F2] = 8'h00;
RAM[16'h14F3] = 8'h00;
RAM[16'h14F4] = 8'h00;
RAM[16'h14F5] = 8'h00;
RAM[16'h14F6] = 8'h00;
RAM[16'h14F7] = 8'h00;
RAM[16'h14F8] = 8'h00;
RAM[16'h14F9] = 8'h00;
RAM[16'h14FA] = 8'h00;
RAM[16'h14FB] = 8'h00;
RAM[16'h14FC] = 8'h00;
RAM[16'h14FD] = 8'h00;
RAM[16'h14FE] = 8'h00;
RAM[16'h14FF] = 8'h00;
RAM[16'h1500] = 8'h00;
RAM[16'h1501] = 8'h00;
RAM[16'h1502] = 8'h00;
RAM[16'h1503] = 8'h00;
RAM[16'h1504] = 8'h00;
RAM[16'h1505] = 8'h00;
RAM[16'h1506] = 8'h00;
RAM[16'h1507] = 8'h00;
RAM[16'h1508] = 8'h00;
RAM[16'h1509] = 8'h00;
RAM[16'h150A] = 8'h00;
RAM[16'h150B] = 8'h00;
RAM[16'h150C] = 8'h00;
RAM[16'h150D] = 8'h00;
RAM[16'h150E] = 8'h00;
RAM[16'h150F] = 8'h00;
RAM[16'h1510] = 8'h00;
RAM[16'h1511] = 8'h00;
RAM[16'h1512] = 8'h00;
RAM[16'h1513] = 8'h00;
RAM[16'h1514] = 8'h00;
RAM[16'h1515] = 8'h00;
RAM[16'h1516] = 8'h00;
RAM[16'h1517] = 8'h00;
RAM[16'h1518] = 8'h00;
RAM[16'h1519] = 8'h00;
RAM[16'h151A] = 8'h00;
RAM[16'h151B] = 8'h00;
RAM[16'h151C] = 8'h00;
RAM[16'h151D] = 8'h00;
RAM[16'h151E] = 8'h00;
RAM[16'h151F] = 8'h00;
RAM[16'h1520] = 8'h00;
RAM[16'h1521] = 8'h00;
RAM[16'h1522] = 8'h00;
RAM[16'h1523] = 8'h00;
RAM[16'h1524] = 8'h00;
RAM[16'h1525] = 8'h00;
RAM[16'h1526] = 8'h00;
RAM[16'h1527] = 8'h00;
RAM[16'h1528] = 8'h00;
RAM[16'h1529] = 8'h00;
RAM[16'h152A] = 8'h00;
RAM[16'h152B] = 8'h00;
RAM[16'h152C] = 8'h00;
RAM[16'h152D] = 8'h00;
RAM[16'h152E] = 8'h00;
RAM[16'h152F] = 8'h00;
RAM[16'h1530] = 8'h00;
RAM[16'h1531] = 8'h00;
RAM[16'h1532] = 8'h00;
RAM[16'h1533] = 8'h00;
RAM[16'h1534] = 8'h00;
RAM[16'h1535] = 8'h00;
RAM[16'h1536] = 8'h00;
RAM[16'h1537] = 8'h00;
RAM[16'h1538] = 8'h00;
RAM[16'h1539] = 8'h00;
RAM[16'h153A] = 8'h00;
RAM[16'h153B] = 8'h00;
RAM[16'h153C] = 8'h00;
RAM[16'h153D] = 8'h00;
RAM[16'h153E] = 8'h00;
RAM[16'h153F] = 8'h00;
RAM[16'h1540] = 8'h00;
RAM[16'h1541] = 8'h00;
RAM[16'h1542] = 8'h00;
RAM[16'h1543] = 8'h00;
RAM[16'h1544] = 8'h00;
RAM[16'h1545] = 8'h00;
RAM[16'h1546] = 8'h00;
RAM[16'h1547] = 8'h00;
RAM[16'h1548] = 8'h00;
RAM[16'h1549] = 8'h00;
RAM[16'h154A] = 8'h00;
RAM[16'h154B] = 8'h00;
RAM[16'h154C] = 8'h00;
RAM[16'h154D] = 8'h00;
RAM[16'h154E] = 8'h00;
RAM[16'h154F] = 8'h00;
RAM[16'h1550] = 8'h00;
RAM[16'h1551] = 8'h00;
RAM[16'h1552] = 8'h00;
RAM[16'h1553] = 8'h00;
RAM[16'h1554] = 8'h00;
RAM[16'h1555] = 8'h00;
RAM[16'h1556] = 8'h00;
RAM[16'h1557] = 8'h00;
RAM[16'h1558] = 8'h00;
RAM[16'h1559] = 8'h00;
RAM[16'h155A] = 8'h00;
RAM[16'h155B] = 8'h00;
RAM[16'h155C] = 8'h00;
RAM[16'h155D] = 8'h00;
RAM[16'h155E] = 8'h00;
RAM[16'h155F] = 8'h00;
RAM[16'h1560] = 8'h00;
RAM[16'h1561] = 8'h00;
RAM[16'h1562] = 8'h00;
RAM[16'h1563] = 8'h00;
RAM[16'h1564] = 8'h00;
RAM[16'h1565] = 8'h00;
RAM[16'h1566] = 8'h00;
RAM[16'h1567] = 8'h00;
RAM[16'h1568] = 8'h00;
RAM[16'h1569] = 8'h00;
RAM[16'h156A] = 8'h00;
RAM[16'h156B] = 8'h00;
RAM[16'h156C] = 8'h00;
RAM[16'h156D] = 8'h00;
RAM[16'h156E] = 8'h00;
RAM[16'h156F] = 8'h00;
RAM[16'h1570] = 8'h00;
RAM[16'h1571] = 8'h00;
RAM[16'h1572] = 8'h00;
RAM[16'h1573] = 8'h00;
RAM[16'h1574] = 8'h00;
RAM[16'h1575] = 8'h00;
RAM[16'h1576] = 8'h00;
RAM[16'h1577] = 8'h00;
RAM[16'h1578] = 8'h00;
RAM[16'h1579] = 8'h00;
RAM[16'h157A] = 8'h00;
RAM[16'h157B] = 8'h00;
RAM[16'h157C] = 8'h00;
RAM[16'h157D] = 8'h00;
RAM[16'h157E] = 8'h00;
RAM[16'h157F] = 8'h00;
RAM[16'h1580] = 8'h00;
RAM[16'h1581] = 8'h00;
RAM[16'h1582] = 8'h00;
RAM[16'h1583] = 8'h00;
RAM[16'h1584] = 8'h00;
RAM[16'h1585] = 8'h00;
RAM[16'h1586] = 8'h00;
RAM[16'h1587] = 8'h00;
RAM[16'h1588] = 8'h00;
RAM[16'h1589] = 8'h00;
RAM[16'h158A] = 8'h00;
RAM[16'h158B] = 8'h00;
RAM[16'h158C] = 8'h00;
RAM[16'h158D] = 8'h00;
RAM[16'h158E] = 8'h00;
RAM[16'h158F] = 8'h00;
RAM[16'h1590] = 8'h00;
RAM[16'h1591] = 8'h00;
RAM[16'h1592] = 8'h00;
RAM[16'h1593] = 8'h00;
RAM[16'h1594] = 8'h00;
RAM[16'h1595] = 8'h00;
RAM[16'h1596] = 8'h00;
RAM[16'h1597] = 8'h00;
RAM[16'h1598] = 8'h00;
RAM[16'h1599] = 8'h00;
RAM[16'h159A] = 8'h00;
RAM[16'h159B] = 8'h00;
RAM[16'h159C] = 8'h00;
RAM[16'h159D] = 8'h00;
RAM[16'h159E] = 8'h00;
RAM[16'h159F] = 8'h00;
RAM[16'h15A0] = 8'h00;
RAM[16'h15A1] = 8'h00;
RAM[16'h15A2] = 8'h00;
RAM[16'h15A3] = 8'h00;
RAM[16'h15A4] = 8'h00;
RAM[16'h15A5] = 8'h00;
RAM[16'h15A6] = 8'h00;
RAM[16'h15A7] = 8'h00;
RAM[16'h15A8] = 8'h00;
RAM[16'h15A9] = 8'h00;
RAM[16'h15AA] = 8'h00;
RAM[16'h15AB] = 8'h00;
RAM[16'h15AC] = 8'h00;
RAM[16'h15AD] = 8'h00;
RAM[16'h15AE] = 8'h00;
RAM[16'h15AF] = 8'h00;
RAM[16'h15B0] = 8'h00;
RAM[16'h15B1] = 8'h00;
RAM[16'h15B2] = 8'h00;
RAM[16'h15B3] = 8'h00;
RAM[16'h15B4] = 8'h00;
RAM[16'h15B5] = 8'h00;
RAM[16'h15B6] = 8'h00;
RAM[16'h15B7] = 8'h00;
RAM[16'h15B8] = 8'h00;
RAM[16'h15B9] = 8'h00;
RAM[16'h15BA] = 8'h00;
RAM[16'h15BB] = 8'h00;
RAM[16'h15BC] = 8'h00;
RAM[16'h15BD] = 8'h00;
RAM[16'h15BE] = 8'h00;
RAM[16'h15BF] = 8'h00;
RAM[16'h15C0] = 8'h00;
RAM[16'h15C1] = 8'h00;
RAM[16'h15C2] = 8'h00;
RAM[16'h15C3] = 8'h00;
RAM[16'h15C4] = 8'h00;
RAM[16'h15C5] = 8'h00;
RAM[16'h15C6] = 8'h00;
RAM[16'h15C7] = 8'h00;
RAM[16'h15C8] = 8'h00;
RAM[16'h15C9] = 8'h00;
RAM[16'h15CA] = 8'h00;
RAM[16'h15CB] = 8'h00;
RAM[16'h15CC] = 8'h00;
RAM[16'h15CD] = 8'h00;
RAM[16'h15CE] = 8'h00;
RAM[16'h15CF] = 8'h00;
RAM[16'h15D0] = 8'h00;
RAM[16'h15D1] = 8'h00;
RAM[16'h15D2] = 8'h00;
RAM[16'h15D3] = 8'h00;
RAM[16'h15D4] = 8'h00;
RAM[16'h15D5] = 8'h00;
RAM[16'h15D6] = 8'h00;
RAM[16'h15D7] = 8'h00;
RAM[16'h15D8] = 8'h00;
RAM[16'h15D9] = 8'h00;
RAM[16'h15DA] = 8'h00;
RAM[16'h15DB] = 8'h00;
RAM[16'h15DC] = 8'h00;
RAM[16'h15DD] = 8'h00;
RAM[16'h15DE] = 8'h00;
RAM[16'h15DF] = 8'h00;
RAM[16'h15E0] = 8'h00;
RAM[16'h15E1] = 8'h00;
RAM[16'h15E2] = 8'h00;
RAM[16'h15E3] = 8'h00;
RAM[16'h15E4] = 8'h00;
RAM[16'h15E5] = 8'h00;
RAM[16'h15E6] = 8'h00;
RAM[16'h15E7] = 8'h00;
RAM[16'h15E8] = 8'h00;
RAM[16'h15E9] = 8'h00;
RAM[16'h15EA] = 8'h00;
RAM[16'h15EB] = 8'h00;
RAM[16'h15EC] = 8'h00;
RAM[16'h15ED] = 8'h00;
RAM[16'h15EE] = 8'h00;
RAM[16'h15EF] = 8'h00;
RAM[16'h15F0] = 8'h00;
RAM[16'h15F1] = 8'h00;
RAM[16'h15F2] = 8'h00;
RAM[16'h15F3] = 8'h00;
RAM[16'h15F4] = 8'h00;
RAM[16'h15F5] = 8'h00;
RAM[16'h15F6] = 8'h00;
RAM[16'h15F7] = 8'h00;
RAM[16'h15F8] = 8'h00;
RAM[16'h15F9] = 8'h00;
RAM[16'h15FA] = 8'h00;
RAM[16'h15FB] = 8'h00;
RAM[16'h15FC] = 8'h00;
RAM[16'h15FD] = 8'h00;
RAM[16'h15FE] = 8'h00;
RAM[16'h15FF] = 8'h00;
RAM[16'h1600] = 8'h00;
RAM[16'h1601] = 8'h00;
RAM[16'h1602] = 8'h00;
RAM[16'h1603] = 8'h00;
RAM[16'h1604] = 8'h00;
RAM[16'h1605] = 8'h00;
RAM[16'h1606] = 8'h00;
RAM[16'h1607] = 8'h00;
RAM[16'h1608] = 8'h00;
RAM[16'h1609] = 8'h00;
RAM[16'h160A] = 8'h00;
RAM[16'h160B] = 8'h00;
RAM[16'h160C] = 8'h00;
RAM[16'h160D] = 8'h00;
RAM[16'h160E] = 8'h00;
RAM[16'h160F] = 8'h00;
RAM[16'h1610] = 8'h00;
RAM[16'h1611] = 8'h00;
RAM[16'h1612] = 8'h00;
RAM[16'h1613] = 8'h00;
RAM[16'h1614] = 8'h00;
RAM[16'h1615] = 8'h00;
RAM[16'h1616] = 8'h00;
RAM[16'h1617] = 8'h00;
RAM[16'h1618] = 8'h00;
RAM[16'h1619] = 8'h00;
RAM[16'h161A] = 8'h00;
RAM[16'h161B] = 8'h00;
RAM[16'h161C] = 8'h00;
RAM[16'h161D] = 8'h00;
RAM[16'h161E] = 8'h00;
RAM[16'h161F] = 8'h00;
RAM[16'h1620] = 8'h00;
RAM[16'h1621] = 8'h00;
RAM[16'h1622] = 8'h00;
RAM[16'h1623] = 8'h00;
RAM[16'h1624] = 8'h00;
RAM[16'h1625] = 8'h00;
RAM[16'h1626] = 8'h00;
RAM[16'h1627] = 8'h00;
RAM[16'h1628] = 8'h00;
RAM[16'h1629] = 8'h00;
RAM[16'h162A] = 8'h00;
RAM[16'h162B] = 8'h00;
RAM[16'h162C] = 8'h00;
RAM[16'h162D] = 8'h00;
RAM[16'h162E] = 8'h00;
RAM[16'h162F] = 8'h00;
RAM[16'h1630] = 8'h00;
RAM[16'h1631] = 8'h00;
RAM[16'h1632] = 8'h00;
RAM[16'h1633] = 8'h00;
RAM[16'h1634] = 8'h00;
RAM[16'h1635] = 8'h00;
RAM[16'h1636] = 8'h00;
RAM[16'h1637] = 8'h00;
RAM[16'h1638] = 8'h00;
RAM[16'h1639] = 8'h00;
RAM[16'h163A] = 8'h00;
RAM[16'h163B] = 8'h00;
RAM[16'h163C] = 8'h00;
RAM[16'h163D] = 8'h00;
RAM[16'h163E] = 8'h00;
RAM[16'h163F] = 8'h00;
RAM[16'h1640] = 8'h00;
RAM[16'h1641] = 8'h00;
RAM[16'h1642] = 8'h00;
RAM[16'h1643] = 8'h00;
RAM[16'h1644] = 8'h00;
RAM[16'h1645] = 8'h00;
RAM[16'h1646] = 8'h00;
RAM[16'h1647] = 8'h00;
RAM[16'h1648] = 8'h00;
RAM[16'h1649] = 8'h00;
RAM[16'h164A] = 8'h00;
RAM[16'h164B] = 8'h00;
RAM[16'h164C] = 8'h00;
RAM[16'h164D] = 8'h00;
RAM[16'h164E] = 8'h00;
RAM[16'h164F] = 8'h00;
RAM[16'h1650] = 8'h00;
RAM[16'h1651] = 8'h00;
RAM[16'h1652] = 8'h00;
RAM[16'h1653] = 8'h00;
RAM[16'h1654] = 8'h00;
RAM[16'h1655] = 8'h00;
RAM[16'h1656] = 8'h00;
RAM[16'h1657] = 8'h00;
RAM[16'h1658] = 8'h00;
RAM[16'h1659] = 8'h00;
RAM[16'h165A] = 8'h00;
RAM[16'h165B] = 8'h00;
RAM[16'h165C] = 8'h00;
RAM[16'h165D] = 8'h00;
RAM[16'h165E] = 8'h00;
RAM[16'h165F] = 8'h00;
RAM[16'h1660] = 8'h00;
RAM[16'h1661] = 8'h00;
RAM[16'h1662] = 8'h00;
RAM[16'h1663] = 8'h00;
RAM[16'h1664] = 8'h00;
RAM[16'h1665] = 8'h00;
RAM[16'h1666] = 8'h00;
RAM[16'h1667] = 8'h00;
RAM[16'h1668] = 8'h00;
RAM[16'h1669] = 8'h00;
RAM[16'h166A] = 8'h00;
RAM[16'h166B] = 8'h00;
RAM[16'h166C] = 8'h00;
RAM[16'h166D] = 8'h00;
RAM[16'h166E] = 8'h00;
RAM[16'h166F] = 8'h00;
RAM[16'h1670] = 8'h00;
RAM[16'h1671] = 8'h00;
RAM[16'h1672] = 8'h00;
RAM[16'h1673] = 8'h00;
RAM[16'h1674] = 8'h00;
RAM[16'h1675] = 8'h00;
RAM[16'h1676] = 8'h00;
RAM[16'h1677] = 8'h00;
RAM[16'h1678] = 8'h00;
RAM[16'h1679] = 8'h00;
RAM[16'h167A] = 8'h00;
RAM[16'h167B] = 8'h00;
RAM[16'h167C] = 8'h00;
RAM[16'h167D] = 8'h00;
RAM[16'h167E] = 8'h00;
RAM[16'h167F] = 8'h00;
RAM[16'h1680] = 8'h00;
RAM[16'h1681] = 8'h00;
RAM[16'h1682] = 8'h00;
RAM[16'h1683] = 8'h00;
RAM[16'h1684] = 8'h00;
RAM[16'h1685] = 8'h00;
RAM[16'h1686] = 8'h00;
RAM[16'h1687] = 8'h00;
RAM[16'h1688] = 8'h00;
RAM[16'h1689] = 8'h00;
RAM[16'h168A] = 8'h00;
RAM[16'h168B] = 8'h00;
RAM[16'h168C] = 8'h00;
RAM[16'h168D] = 8'h00;
RAM[16'h168E] = 8'h00;
RAM[16'h168F] = 8'h00;
RAM[16'h1690] = 8'h00;
RAM[16'h1691] = 8'h00;
RAM[16'h1692] = 8'h00;
RAM[16'h1693] = 8'h00;
RAM[16'h1694] = 8'h00;
RAM[16'h1695] = 8'h00;
RAM[16'h1696] = 8'h00;
RAM[16'h1697] = 8'h00;
RAM[16'h1698] = 8'h00;
RAM[16'h1699] = 8'h00;
RAM[16'h169A] = 8'h00;
RAM[16'h169B] = 8'h00;
RAM[16'h169C] = 8'h00;
RAM[16'h169D] = 8'h00;
RAM[16'h169E] = 8'h00;
RAM[16'h169F] = 8'h00;
RAM[16'h16A0] = 8'h00;
RAM[16'h16A1] = 8'h00;
RAM[16'h16A2] = 8'h00;
RAM[16'h16A3] = 8'h00;
RAM[16'h16A4] = 8'h00;
RAM[16'h16A5] = 8'h00;
RAM[16'h16A6] = 8'h00;
RAM[16'h16A7] = 8'h00;
RAM[16'h16A8] = 8'h00;
RAM[16'h16A9] = 8'h00;
RAM[16'h16AA] = 8'h00;
RAM[16'h16AB] = 8'h00;
RAM[16'h16AC] = 8'h00;
RAM[16'h16AD] = 8'h00;
RAM[16'h16AE] = 8'h00;
RAM[16'h16AF] = 8'h00;
RAM[16'h16B0] = 8'h00;
RAM[16'h16B1] = 8'h00;
RAM[16'h16B2] = 8'h00;
RAM[16'h16B3] = 8'h00;
RAM[16'h16B4] = 8'h00;
RAM[16'h16B5] = 8'h00;
RAM[16'h16B6] = 8'h00;
RAM[16'h16B7] = 8'h00;
RAM[16'h16B8] = 8'h00;
RAM[16'h16B9] = 8'h00;
RAM[16'h16BA] = 8'h00;
RAM[16'h16BB] = 8'h00;
RAM[16'h16BC] = 8'h00;
RAM[16'h16BD] = 8'h00;
RAM[16'h16BE] = 8'h00;
RAM[16'h16BF] = 8'h00;
RAM[16'h16C0] = 8'h00;
RAM[16'h16C1] = 8'h00;
RAM[16'h16C2] = 8'h00;
RAM[16'h16C3] = 8'h00;
RAM[16'h16C4] = 8'h00;
RAM[16'h16C5] = 8'h00;
RAM[16'h16C6] = 8'h00;
RAM[16'h16C7] = 8'h00;
RAM[16'h16C8] = 8'h00;
RAM[16'h16C9] = 8'h00;
RAM[16'h16CA] = 8'h00;
RAM[16'h16CB] = 8'h00;
RAM[16'h16CC] = 8'h00;
RAM[16'h16CD] = 8'h00;
RAM[16'h16CE] = 8'h00;
RAM[16'h16CF] = 8'h00;
RAM[16'h16D0] = 8'h00;
RAM[16'h16D1] = 8'h00;
RAM[16'h16D2] = 8'h00;
RAM[16'h16D3] = 8'h00;
RAM[16'h16D4] = 8'h00;
RAM[16'h16D5] = 8'h00;
RAM[16'h16D6] = 8'h00;
RAM[16'h16D7] = 8'h00;
RAM[16'h16D8] = 8'h00;
RAM[16'h16D9] = 8'h00;
RAM[16'h16DA] = 8'h00;
RAM[16'h16DB] = 8'h00;
RAM[16'h16DC] = 8'h00;
RAM[16'h16DD] = 8'h00;
RAM[16'h16DE] = 8'h00;
RAM[16'h16DF] = 8'h00;
RAM[16'h16E0] = 8'h00;
RAM[16'h16E1] = 8'h00;
RAM[16'h16E2] = 8'h00;
RAM[16'h16E3] = 8'h00;
RAM[16'h16E4] = 8'h00;
RAM[16'h16E5] = 8'h00;
RAM[16'h16E6] = 8'h00;
RAM[16'h16E7] = 8'h00;
RAM[16'h16E8] = 8'h00;
RAM[16'h16E9] = 8'h00;
RAM[16'h16EA] = 8'h00;
RAM[16'h16EB] = 8'h00;
RAM[16'h16EC] = 8'h00;
RAM[16'h16ED] = 8'h00;
RAM[16'h16EE] = 8'h00;
RAM[16'h16EF] = 8'h00;
RAM[16'h16F0] = 8'h00;
RAM[16'h16F1] = 8'h00;
RAM[16'h16F2] = 8'h00;
RAM[16'h16F3] = 8'h00;
RAM[16'h16F4] = 8'h00;
RAM[16'h16F5] = 8'h00;
RAM[16'h16F6] = 8'h00;
RAM[16'h16F7] = 8'h00;
RAM[16'h16F8] = 8'h00;
RAM[16'h16F9] = 8'h00;
RAM[16'h16FA] = 8'h00;
RAM[16'h16FB] = 8'h00;
RAM[16'h16FC] = 8'h00;
RAM[16'h16FD] = 8'h00;
RAM[16'h16FE] = 8'h00;
RAM[16'h16FF] = 8'h00;
RAM[16'h1700] = 8'h00;
RAM[16'h1701] = 8'h00;
RAM[16'h1702] = 8'h00;
RAM[16'h1703] = 8'h00;
RAM[16'h1704] = 8'h00;
RAM[16'h1705] = 8'h00;
RAM[16'h1706] = 8'h00;
RAM[16'h1707] = 8'h00;
RAM[16'h1708] = 8'h00;
RAM[16'h1709] = 8'h00;
RAM[16'h170A] = 8'h00;
RAM[16'h170B] = 8'h00;
RAM[16'h170C] = 8'h00;
RAM[16'h170D] = 8'h00;
RAM[16'h170E] = 8'h00;
RAM[16'h170F] = 8'h00;
RAM[16'h1710] = 8'h00;
RAM[16'h1711] = 8'h00;
RAM[16'h1712] = 8'h00;
RAM[16'h1713] = 8'h00;
RAM[16'h1714] = 8'h00;
RAM[16'h1715] = 8'h00;
RAM[16'h1716] = 8'h00;
RAM[16'h1717] = 8'h00;
RAM[16'h1718] = 8'h00;
RAM[16'h1719] = 8'h00;
RAM[16'h171A] = 8'h00;
RAM[16'h171B] = 8'h00;
RAM[16'h171C] = 8'h00;
RAM[16'h171D] = 8'h00;
RAM[16'h171E] = 8'h00;
RAM[16'h171F] = 8'h00;
RAM[16'h1720] = 8'h00;
RAM[16'h1721] = 8'h00;
RAM[16'h1722] = 8'h00;
RAM[16'h1723] = 8'h00;
RAM[16'h1724] = 8'h00;
RAM[16'h1725] = 8'h00;
RAM[16'h1726] = 8'h00;
RAM[16'h1727] = 8'h00;
RAM[16'h1728] = 8'h00;
RAM[16'h1729] = 8'h00;
RAM[16'h172A] = 8'h00;
RAM[16'h172B] = 8'h00;
RAM[16'h172C] = 8'h00;
RAM[16'h172D] = 8'h00;
RAM[16'h172E] = 8'h00;
RAM[16'h172F] = 8'h00;
RAM[16'h1730] = 8'h00;
RAM[16'h1731] = 8'h00;
RAM[16'h1732] = 8'h00;
RAM[16'h1733] = 8'h00;
RAM[16'h1734] = 8'h00;
RAM[16'h1735] = 8'h00;
RAM[16'h1736] = 8'h00;
RAM[16'h1737] = 8'h00;
RAM[16'h1738] = 8'h00;
RAM[16'h1739] = 8'h00;
RAM[16'h173A] = 8'h00;
RAM[16'h173B] = 8'h00;
RAM[16'h173C] = 8'h00;
RAM[16'h173D] = 8'h00;
RAM[16'h173E] = 8'h00;
RAM[16'h173F] = 8'h00;
RAM[16'h1740] = 8'h00;
RAM[16'h1741] = 8'h00;
RAM[16'h1742] = 8'h00;
RAM[16'h1743] = 8'h00;
RAM[16'h1744] = 8'h00;
RAM[16'h1745] = 8'h00;
RAM[16'h1746] = 8'h00;
RAM[16'h1747] = 8'h00;
RAM[16'h1748] = 8'h00;
RAM[16'h1749] = 8'h00;
RAM[16'h174A] = 8'h00;
RAM[16'h174B] = 8'h00;
RAM[16'h174C] = 8'h00;
RAM[16'h174D] = 8'h00;
RAM[16'h174E] = 8'h00;
RAM[16'h174F] = 8'h00;
RAM[16'h1750] = 8'h00;
RAM[16'h1751] = 8'h00;
RAM[16'h1752] = 8'h00;
RAM[16'h1753] = 8'h00;
RAM[16'h1754] = 8'h00;
RAM[16'h1755] = 8'h00;
RAM[16'h1756] = 8'h00;
RAM[16'h1757] = 8'h00;
RAM[16'h1758] = 8'h00;
RAM[16'h1759] = 8'h00;
RAM[16'h175A] = 8'h00;
RAM[16'h175B] = 8'h00;
RAM[16'h175C] = 8'h00;
RAM[16'h175D] = 8'h00;
RAM[16'h175E] = 8'h00;
RAM[16'h175F] = 8'h00;
RAM[16'h1760] = 8'h00;
RAM[16'h1761] = 8'h00;
RAM[16'h1762] = 8'h00;
RAM[16'h1763] = 8'h00;
RAM[16'h1764] = 8'h00;
RAM[16'h1765] = 8'h00;
RAM[16'h1766] = 8'h00;
RAM[16'h1767] = 8'h00;
RAM[16'h1768] = 8'h00;
RAM[16'h1769] = 8'h00;
RAM[16'h176A] = 8'h00;
RAM[16'h176B] = 8'h00;
RAM[16'h176C] = 8'h00;
RAM[16'h176D] = 8'h00;
RAM[16'h176E] = 8'h00;
RAM[16'h176F] = 8'h00;
RAM[16'h1770] = 8'h00;
RAM[16'h1771] = 8'h00;
RAM[16'h1772] = 8'h00;
RAM[16'h1773] = 8'h00;
RAM[16'h1774] = 8'h00;
RAM[16'h1775] = 8'h00;
RAM[16'h1776] = 8'h00;
RAM[16'h1777] = 8'h00;
RAM[16'h1778] = 8'h00;
RAM[16'h1779] = 8'h00;
RAM[16'h177A] = 8'h00;
RAM[16'h177B] = 8'h00;
RAM[16'h177C] = 8'h00;
RAM[16'h177D] = 8'h00;
RAM[16'h177E] = 8'h00;
RAM[16'h177F] = 8'h00;
RAM[16'h1780] = 8'h00;
RAM[16'h1781] = 8'h00;
RAM[16'h1782] = 8'h00;
RAM[16'h1783] = 8'h00;
RAM[16'h1784] = 8'h00;
RAM[16'h1785] = 8'h00;
RAM[16'h1786] = 8'h00;
RAM[16'h1787] = 8'h00;
RAM[16'h1788] = 8'h00;
RAM[16'h1789] = 8'h00;
RAM[16'h178A] = 8'h00;
RAM[16'h178B] = 8'h00;
RAM[16'h178C] = 8'h00;
RAM[16'h178D] = 8'h00;
RAM[16'h178E] = 8'h00;
RAM[16'h178F] = 8'h00;
RAM[16'h1790] = 8'h00;
RAM[16'h1791] = 8'h00;
RAM[16'h1792] = 8'h00;
RAM[16'h1793] = 8'h00;
RAM[16'h1794] = 8'h00;
RAM[16'h1795] = 8'h00;
RAM[16'h1796] = 8'h00;
RAM[16'h1797] = 8'h00;
RAM[16'h1798] = 8'h00;
RAM[16'h1799] = 8'h00;
RAM[16'h179A] = 8'h00;
RAM[16'h179B] = 8'h00;
RAM[16'h179C] = 8'h00;
RAM[16'h179D] = 8'h00;
RAM[16'h179E] = 8'h00;
RAM[16'h179F] = 8'h00;
RAM[16'h17A0] = 8'h00;
RAM[16'h17A1] = 8'h00;
RAM[16'h17A2] = 8'h00;
RAM[16'h17A3] = 8'h00;
RAM[16'h17A4] = 8'h00;
RAM[16'h17A5] = 8'h00;
RAM[16'h17A6] = 8'h00;
RAM[16'h17A7] = 8'h00;
RAM[16'h17A8] = 8'h00;
RAM[16'h17A9] = 8'h00;
RAM[16'h17AA] = 8'h00;
RAM[16'h17AB] = 8'h00;
RAM[16'h17AC] = 8'h00;
RAM[16'h17AD] = 8'h00;
RAM[16'h17AE] = 8'h00;
RAM[16'h17AF] = 8'h00;
RAM[16'h17B0] = 8'h00;
RAM[16'h17B1] = 8'h00;
RAM[16'h17B2] = 8'h00;
RAM[16'h17B3] = 8'h00;
RAM[16'h17B4] = 8'h00;
RAM[16'h17B5] = 8'h00;
RAM[16'h17B6] = 8'h00;
RAM[16'h17B7] = 8'h00;
RAM[16'h17B8] = 8'h00;
RAM[16'h17B9] = 8'h00;
RAM[16'h17BA] = 8'h00;
RAM[16'h17BB] = 8'h00;
RAM[16'h17BC] = 8'h00;
RAM[16'h17BD] = 8'h00;
RAM[16'h17BE] = 8'h00;
RAM[16'h17BF] = 8'h00;
RAM[16'h17C0] = 8'h00;
RAM[16'h17C1] = 8'h00;
RAM[16'h17C2] = 8'h00;
RAM[16'h17C3] = 8'h00;
RAM[16'h17C4] = 8'h00;
RAM[16'h17C5] = 8'h00;
RAM[16'h17C6] = 8'h00;
RAM[16'h17C7] = 8'h00;
RAM[16'h17C8] = 8'h00;
RAM[16'h17C9] = 8'h00;
RAM[16'h17CA] = 8'h00;
RAM[16'h17CB] = 8'h00;
RAM[16'h17CC] = 8'h00;
RAM[16'h17CD] = 8'h00;
RAM[16'h17CE] = 8'h00;
RAM[16'h17CF] = 8'h00;
RAM[16'h17D0] = 8'h00;
RAM[16'h17D1] = 8'h00;
RAM[16'h17D2] = 8'h00;
RAM[16'h17D3] = 8'h00;
RAM[16'h17D4] = 8'h00;
RAM[16'h17D5] = 8'h00;
RAM[16'h17D6] = 8'h00;
RAM[16'h17D7] = 8'h00;
RAM[16'h17D8] = 8'h00;
RAM[16'h17D9] = 8'h00;
RAM[16'h17DA] = 8'h00;
RAM[16'h17DB] = 8'h00;
RAM[16'h17DC] = 8'h00;
RAM[16'h17DD] = 8'h00;
RAM[16'h17DE] = 8'h00;
RAM[16'h17DF] = 8'h00;
RAM[16'h17E0] = 8'h00;
RAM[16'h17E1] = 8'h00;
RAM[16'h17E2] = 8'h00;
RAM[16'h17E3] = 8'h00;
RAM[16'h17E4] = 8'h00;
RAM[16'h17E5] = 8'h00;
RAM[16'h17E6] = 8'h00;
RAM[16'h17E7] = 8'h00;
RAM[16'h17E8] = 8'h00;
RAM[16'h17E9] = 8'h00;
RAM[16'h17EA] = 8'h00;
RAM[16'h17EB] = 8'h00;
RAM[16'h17EC] = 8'h00;
RAM[16'h17ED] = 8'h00;
RAM[16'h17EE] = 8'h00;
RAM[16'h17EF] = 8'h00;
RAM[16'h17F0] = 8'h00;
RAM[16'h17F1] = 8'h00;
RAM[16'h17F2] = 8'h00;
RAM[16'h17F3] = 8'h00;
RAM[16'h17F4] = 8'h00;
RAM[16'h17F5] = 8'h00;
RAM[16'h17F6] = 8'h00;
RAM[16'h17F7] = 8'h00;
RAM[16'h17F8] = 8'h00;
RAM[16'h17F9] = 8'h00;
RAM[16'h17FA] = 8'h00;
RAM[16'h17FB] = 8'h00;
RAM[16'h17FC] = 8'h00;
RAM[16'h17FD] = 8'h00;
RAM[16'h17FE] = 8'h00;
RAM[16'h17FF] = 8'h00;
RAM[16'h1800] = 8'h00;
RAM[16'h1801] = 8'h00;
RAM[16'h1802] = 8'h00;
RAM[16'h1803] = 8'h00;
RAM[16'h1804] = 8'h00;
RAM[16'h1805] = 8'h00;
RAM[16'h1806] = 8'h00;
RAM[16'h1807] = 8'h00;
RAM[16'h1808] = 8'h00;
RAM[16'h1809] = 8'h00;
RAM[16'h180A] = 8'h00;
RAM[16'h180B] = 8'h00;
RAM[16'h180C] = 8'h00;
RAM[16'h180D] = 8'h00;
RAM[16'h180E] = 8'h00;
RAM[16'h180F] = 8'h00;
RAM[16'h1810] = 8'h00;
RAM[16'h1811] = 8'h00;
RAM[16'h1812] = 8'h00;
RAM[16'h1813] = 8'h00;
RAM[16'h1814] = 8'h00;
RAM[16'h1815] = 8'h00;
RAM[16'h1816] = 8'h00;
RAM[16'h1817] = 8'h00;
RAM[16'h1818] = 8'h00;
RAM[16'h1819] = 8'h00;
RAM[16'h181A] = 8'h00;
RAM[16'h181B] = 8'h00;
RAM[16'h181C] = 8'h00;
RAM[16'h181D] = 8'h00;
RAM[16'h181E] = 8'h00;
RAM[16'h181F] = 8'h00;
RAM[16'h1820] = 8'h00;
RAM[16'h1821] = 8'h00;
RAM[16'h1822] = 8'h00;
RAM[16'h1823] = 8'h00;
RAM[16'h1824] = 8'h00;
RAM[16'h1825] = 8'h00;
RAM[16'h1826] = 8'h00;
RAM[16'h1827] = 8'h00;
RAM[16'h1828] = 8'h00;
RAM[16'h1829] = 8'h00;
RAM[16'h182A] = 8'h00;
RAM[16'h182B] = 8'h00;
RAM[16'h182C] = 8'h00;
RAM[16'h182D] = 8'h00;
RAM[16'h182E] = 8'h00;
RAM[16'h182F] = 8'h00;
RAM[16'h1830] = 8'h00;
RAM[16'h1831] = 8'h00;
RAM[16'h1832] = 8'h00;
RAM[16'h1833] = 8'h00;
RAM[16'h1834] = 8'h00;
RAM[16'h1835] = 8'h00;
RAM[16'h1836] = 8'h00;
RAM[16'h1837] = 8'h00;
RAM[16'h1838] = 8'h00;
RAM[16'h1839] = 8'h00;
RAM[16'h183A] = 8'h00;
RAM[16'h183B] = 8'h00;
RAM[16'h183C] = 8'h00;
RAM[16'h183D] = 8'h00;
RAM[16'h183E] = 8'h00;
RAM[16'h183F] = 8'h00;
RAM[16'h1840] = 8'h00;
RAM[16'h1841] = 8'h00;
RAM[16'h1842] = 8'h00;
RAM[16'h1843] = 8'h00;
RAM[16'h1844] = 8'h00;
RAM[16'h1845] = 8'h00;
RAM[16'h1846] = 8'h00;
RAM[16'h1847] = 8'h00;
RAM[16'h1848] = 8'h00;
RAM[16'h1849] = 8'h00;
RAM[16'h184A] = 8'h00;
RAM[16'h184B] = 8'h00;
RAM[16'h184C] = 8'h00;
RAM[16'h184D] = 8'h00;
RAM[16'h184E] = 8'h00;
RAM[16'h184F] = 8'h00;
RAM[16'h1850] = 8'h00;
RAM[16'h1851] = 8'h00;
RAM[16'h1852] = 8'h00;
RAM[16'h1853] = 8'h00;
RAM[16'h1854] = 8'h00;
RAM[16'h1855] = 8'h00;
RAM[16'h1856] = 8'h00;
RAM[16'h1857] = 8'h00;
RAM[16'h1858] = 8'h00;
RAM[16'h1859] = 8'h00;
RAM[16'h185A] = 8'h00;
RAM[16'h185B] = 8'h00;
RAM[16'h185C] = 8'h00;
RAM[16'h185D] = 8'h00;
RAM[16'h185E] = 8'h00;
RAM[16'h185F] = 8'h00;
RAM[16'h1860] = 8'h00;
RAM[16'h1861] = 8'h00;
RAM[16'h1862] = 8'h00;
RAM[16'h1863] = 8'h00;
RAM[16'h1864] = 8'h00;
RAM[16'h1865] = 8'h00;
RAM[16'h1866] = 8'h00;
RAM[16'h1867] = 8'h00;
RAM[16'h1868] = 8'h00;
RAM[16'h1869] = 8'h00;
RAM[16'h186A] = 8'h00;
RAM[16'h186B] = 8'h00;
RAM[16'h186C] = 8'h00;
RAM[16'h186D] = 8'h00;
RAM[16'h186E] = 8'h00;
RAM[16'h186F] = 8'h00;
RAM[16'h1870] = 8'h00;
RAM[16'h1871] = 8'h00;
RAM[16'h1872] = 8'h00;
RAM[16'h1873] = 8'h00;
RAM[16'h1874] = 8'h00;
RAM[16'h1875] = 8'h00;
RAM[16'h1876] = 8'h00;
RAM[16'h1877] = 8'h00;
RAM[16'h1878] = 8'h00;
RAM[16'h1879] = 8'h00;
RAM[16'h187A] = 8'h00;
RAM[16'h187B] = 8'h00;
RAM[16'h187C] = 8'h00;
RAM[16'h187D] = 8'h00;
RAM[16'h187E] = 8'h00;
RAM[16'h187F] = 8'h00;
RAM[16'h1880] = 8'h00;
RAM[16'h1881] = 8'h00;
RAM[16'h1882] = 8'h00;
RAM[16'h1883] = 8'h00;
RAM[16'h1884] = 8'h00;
RAM[16'h1885] = 8'h00;
RAM[16'h1886] = 8'h00;
RAM[16'h1887] = 8'h00;
RAM[16'h1888] = 8'h00;
RAM[16'h1889] = 8'h00;
RAM[16'h188A] = 8'h00;
RAM[16'h188B] = 8'h00;
RAM[16'h188C] = 8'h00;
RAM[16'h188D] = 8'h00;
RAM[16'h188E] = 8'h00;
RAM[16'h188F] = 8'h00;
RAM[16'h1890] = 8'h00;
RAM[16'h1891] = 8'h00;
RAM[16'h1892] = 8'h00;
RAM[16'h1893] = 8'h00;
RAM[16'h1894] = 8'h00;
RAM[16'h1895] = 8'h00;
RAM[16'h1896] = 8'h00;
RAM[16'h1897] = 8'h00;
RAM[16'h1898] = 8'h00;
RAM[16'h1899] = 8'h00;
RAM[16'h189A] = 8'h00;
RAM[16'h189B] = 8'h00;
RAM[16'h189C] = 8'h00;
RAM[16'h189D] = 8'h00;
RAM[16'h189E] = 8'h00;
RAM[16'h189F] = 8'h00;
RAM[16'h18A0] = 8'h00;
RAM[16'h18A1] = 8'h00;
RAM[16'h18A2] = 8'h00;
RAM[16'h18A3] = 8'h00;
RAM[16'h18A4] = 8'h00;
RAM[16'h18A5] = 8'h00;
RAM[16'h18A6] = 8'h00;
RAM[16'h18A7] = 8'h00;
RAM[16'h18A8] = 8'h00;
RAM[16'h18A9] = 8'h00;
RAM[16'h18AA] = 8'h00;
RAM[16'h18AB] = 8'h00;
RAM[16'h18AC] = 8'h00;
RAM[16'h18AD] = 8'h00;
RAM[16'h18AE] = 8'h00;
RAM[16'h18AF] = 8'h00;
RAM[16'h18B0] = 8'h00;
RAM[16'h18B1] = 8'h00;
RAM[16'h18B2] = 8'h00;
RAM[16'h18B3] = 8'h00;
RAM[16'h18B4] = 8'h00;
RAM[16'h18B5] = 8'h00;
RAM[16'h18B6] = 8'h00;
RAM[16'h18B7] = 8'h00;
RAM[16'h18B8] = 8'h00;
RAM[16'h18B9] = 8'h00;
RAM[16'h18BA] = 8'h00;
RAM[16'h18BB] = 8'h00;
RAM[16'h18BC] = 8'h00;
RAM[16'h18BD] = 8'h00;
RAM[16'h18BE] = 8'h00;
RAM[16'h18BF] = 8'h00;
RAM[16'h18C0] = 8'h00;
RAM[16'h18C1] = 8'h00;
RAM[16'h18C2] = 8'h00;
RAM[16'h18C3] = 8'h00;
RAM[16'h18C4] = 8'h00;
RAM[16'h18C5] = 8'h00;
RAM[16'h18C6] = 8'h00;
RAM[16'h18C7] = 8'h00;
RAM[16'h18C8] = 8'h00;
RAM[16'h18C9] = 8'h00;
RAM[16'h18CA] = 8'h00;
RAM[16'h18CB] = 8'h00;
RAM[16'h18CC] = 8'h00;
RAM[16'h18CD] = 8'h00;
RAM[16'h18CE] = 8'h00;
RAM[16'h18CF] = 8'h00;
RAM[16'h18D0] = 8'h00;
RAM[16'h18D1] = 8'h00;
RAM[16'h18D2] = 8'h00;
RAM[16'h18D3] = 8'h00;
RAM[16'h18D4] = 8'h00;
RAM[16'h18D5] = 8'h00;
RAM[16'h18D6] = 8'h00;
RAM[16'h18D7] = 8'h00;
RAM[16'h18D8] = 8'h00;
RAM[16'h18D9] = 8'h00;
RAM[16'h18DA] = 8'h00;
RAM[16'h18DB] = 8'h00;
RAM[16'h18DC] = 8'h00;
RAM[16'h18DD] = 8'h00;
RAM[16'h18DE] = 8'h00;
RAM[16'h18DF] = 8'h00;
RAM[16'h18E0] = 8'h00;
RAM[16'h18E1] = 8'h00;
RAM[16'h18E2] = 8'h00;
RAM[16'h18E3] = 8'h00;
RAM[16'h18E4] = 8'h00;
RAM[16'h18E5] = 8'h00;
RAM[16'h18E6] = 8'h00;
RAM[16'h18E7] = 8'h00;
RAM[16'h18E8] = 8'h00;
RAM[16'h18E9] = 8'h00;
RAM[16'h18EA] = 8'h00;
RAM[16'h18EB] = 8'h00;
RAM[16'h18EC] = 8'h00;
RAM[16'h18ED] = 8'h00;
RAM[16'h18EE] = 8'h00;
RAM[16'h18EF] = 8'h00;
RAM[16'h18F0] = 8'h00;
RAM[16'h18F1] = 8'h00;
RAM[16'h18F2] = 8'h00;
RAM[16'h18F3] = 8'h00;
RAM[16'h18F4] = 8'h00;
RAM[16'h18F5] = 8'h00;
RAM[16'h18F6] = 8'h00;
RAM[16'h18F7] = 8'h00;
RAM[16'h18F8] = 8'h00;
RAM[16'h18F9] = 8'h00;
RAM[16'h18FA] = 8'h00;
RAM[16'h18FB] = 8'h00;
RAM[16'h18FC] = 8'h00;
RAM[16'h18FD] = 8'h00;
RAM[16'h18FE] = 8'h00;
RAM[16'h18FF] = 8'h00;
RAM[16'h1900] = 8'h00;
RAM[16'h1901] = 8'h00;
RAM[16'h1902] = 8'h00;
RAM[16'h1903] = 8'h00;
RAM[16'h1904] = 8'h00;
RAM[16'h1905] = 8'h00;
RAM[16'h1906] = 8'h00;
RAM[16'h1907] = 8'h00;
RAM[16'h1908] = 8'h00;
RAM[16'h1909] = 8'h00;
RAM[16'h190A] = 8'h00;
RAM[16'h190B] = 8'h00;
RAM[16'h190C] = 8'h00;
RAM[16'h190D] = 8'h00;
RAM[16'h190E] = 8'h00;
RAM[16'h190F] = 8'h00;
RAM[16'h1910] = 8'h00;
RAM[16'h1911] = 8'h00;
RAM[16'h1912] = 8'h00;
RAM[16'h1913] = 8'h00;
RAM[16'h1914] = 8'h00;
RAM[16'h1915] = 8'h00;
RAM[16'h1916] = 8'h00;
RAM[16'h1917] = 8'h00;
RAM[16'h1918] = 8'h00;
RAM[16'h1919] = 8'h00;
RAM[16'h191A] = 8'h00;
RAM[16'h191B] = 8'h00;
RAM[16'h191C] = 8'h00;
RAM[16'h191D] = 8'h00;
RAM[16'h191E] = 8'h00;
RAM[16'h191F] = 8'h00;
RAM[16'h1920] = 8'h00;
RAM[16'h1921] = 8'h00;
RAM[16'h1922] = 8'h00;
RAM[16'h1923] = 8'h00;
RAM[16'h1924] = 8'h00;
RAM[16'h1925] = 8'h00;
RAM[16'h1926] = 8'h00;
RAM[16'h1927] = 8'h00;
RAM[16'h1928] = 8'h00;
RAM[16'h1929] = 8'h00;
RAM[16'h192A] = 8'h00;
RAM[16'h192B] = 8'h00;
RAM[16'h192C] = 8'h00;
RAM[16'h192D] = 8'h00;
RAM[16'h192E] = 8'h00;
RAM[16'h192F] = 8'h00;
RAM[16'h1930] = 8'h00;
RAM[16'h1931] = 8'h00;
RAM[16'h1932] = 8'h00;
RAM[16'h1933] = 8'h00;
RAM[16'h1934] = 8'h00;
RAM[16'h1935] = 8'h00;
RAM[16'h1936] = 8'h00;
RAM[16'h1937] = 8'h00;
RAM[16'h1938] = 8'h00;
RAM[16'h1939] = 8'h00;
RAM[16'h193A] = 8'h00;
RAM[16'h193B] = 8'h00;
RAM[16'h193C] = 8'h00;
RAM[16'h193D] = 8'h00;
RAM[16'h193E] = 8'h00;
RAM[16'h193F] = 8'h00;
RAM[16'h1940] = 8'h00;
RAM[16'h1941] = 8'h00;
RAM[16'h1942] = 8'h00;
RAM[16'h1943] = 8'h00;
RAM[16'h1944] = 8'h00;
RAM[16'h1945] = 8'h00;
RAM[16'h1946] = 8'h00;
RAM[16'h1947] = 8'h00;
RAM[16'h1948] = 8'h00;
RAM[16'h1949] = 8'h00;
RAM[16'h194A] = 8'h00;
RAM[16'h194B] = 8'h00;
RAM[16'h194C] = 8'h00;
RAM[16'h194D] = 8'h00;
RAM[16'h194E] = 8'h00;
RAM[16'h194F] = 8'h00;
RAM[16'h1950] = 8'h00;
RAM[16'h1951] = 8'h00;
RAM[16'h1952] = 8'h00;
RAM[16'h1953] = 8'h00;
RAM[16'h1954] = 8'h00;
RAM[16'h1955] = 8'h00;
RAM[16'h1956] = 8'h00;
RAM[16'h1957] = 8'h00;
RAM[16'h1958] = 8'h00;
RAM[16'h1959] = 8'h00;
RAM[16'h195A] = 8'h00;
RAM[16'h195B] = 8'h00;
RAM[16'h195C] = 8'h00;
RAM[16'h195D] = 8'h00;
RAM[16'h195E] = 8'h00;
RAM[16'h195F] = 8'h00;
RAM[16'h1960] = 8'h00;
RAM[16'h1961] = 8'h00;
RAM[16'h1962] = 8'h00;
RAM[16'h1963] = 8'h00;
RAM[16'h1964] = 8'h00;
RAM[16'h1965] = 8'h00;
RAM[16'h1966] = 8'h00;
RAM[16'h1967] = 8'h00;
RAM[16'h1968] = 8'h00;
RAM[16'h1969] = 8'h00;
RAM[16'h196A] = 8'h00;
RAM[16'h196B] = 8'h00;
RAM[16'h196C] = 8'h00;
RAM[16'h196D] = 8'h00;
RAM[16'h196E] = 8'h00;
RAM[16'h196F] = 8'h00;
RAM[16'h1970] = 8'h00;
RAM[16'h1971] = 8'h00;
RAM[16'h1972] = 8'h00;
RAM[16'h1973] = 8'h00;
RAM[16'h1974] = 8'h00;
RAM[16'h1975] = 8'h00;
RAM[16'h1976] = 8'h00;
RAM[16'h1977] = 8'h00;
RAM[16'h1978] = 8'h00;
RAM[16'h1979] = 8'h00;
RAM[16'h197A] = 8'h00;
RAM[16'h197B] = 8'h00;
RAM[16'h197C] = 8'h00;
RAM[16'h197D] = 8'h00;
RAM[16'h197E] = 8'h00;
RAM[16'h197F] = 8'h00;
RAM[16'h1980] = 8'h00;
RAM[16'h1981] = 8'h00;
RAM[16'h1982] = 8'h00;
RAM[16'h1983] = 8'h00;
RAM[16'h1984] = 8'h00;
RAM[16'h1985] = 8'h00;
RAM[16'h1986] = 8'h00;
RAM[16'h1987] = 8'h00;
RAM[16'h1988] = 8'h00;
RAM[16'h1989] = 8'h00;
RAM[16'h198A] = 8'h00;
RAM[16'h198B] = 8'h00;
RAM[16'h198C] = 8'h00;
RAM[16'h198D] = 8'h00;
RAM[16'h198E] = 8'h00;
RAM[16'h198F] = 8'h00;
RAM[16'h1990] = 8'h00;
RAM[16'h1991] = 8'h00;
RAM[16'h1992] = 8'h00;
RAM[16'h1993] = 8'h00;
RAM[16'h1994] = 8'h00;
RAM[16'h1995] = 8'h00;
RAM[16'h1996] = 8'h00;
RAM[16'h1997] = 8'h00;
RAM[16'h1998] = 8'h00;
RAM[16'h1999] = 8'h00;
RAM[16'h199A] = 8'h00;
RAM[16'h199B] = 8'h00;
RAM[16'h199C] = 8'h00;
RAM[16'h199D] = 8'h00;
RAM[16'h199E] = 8'h00;
RAM[16'h199F] = 8'h00;
RAM[16'h19A0] = 8'h00;
RAM[16'h19A1] = 8'h00;
RAM[16'h19A2] = 8'h00;
RAM[16'h19A3] = 8'h00;
RAM[16'h19A4] = 8'h00;
RAM[16'h19A5] = 8'h00;
RAM[16'h19A6] = 8'h00;
RAM[16'h19A7] = 8'h00;
RAM[16'h19A8] = 8'h00;
RAM[16'h19A9] = 8'h00;
RAM[16'h19AA] = 8'h00;
RAM[16'h19AB] = 8'h00;
RAM[16'h19AC] = 8'h00;
RAM[16'h19AD] = 8'h00;
RAM[16'h19AE] = 8'h00;
RAM[16'h19AF] = 8'h00;
RAM[16'h19B0] = 8'h00;
RAM[16'h19B1] = 8'h00;
RAM[16'h19B2] = 8'h00;
RAM[16'h19B3] = 8'h00;
RAM[16'h19B4] = 8'h00;
RAM[16'h19B5] = 8'h00;
RAM[16'h19B6] = 8'h00;
RAM[16'h19B7] = 8'h00;
RAM[16'h19B8] = 8'h00;
RAM[16'h19B9] = 8'h00;
RAM[16'h19BA] = 8'h00;
RAM[16'h19BB] = 8'h00;
RAM[16'h19BC] = 8'h00;
RAM[16'h19BD] = 8'h00;
RAM[16'h19BE] = 8'h00;
RAM[16'h19BF] = 8'h00;
RAM[16'h19C0] = 8'h00;
RAM[16'h19C1] = 8'h00;
RAM[16'h19C2] = 8'h00;
RAM[16'h19C3] = 8'h00;
RAM[16'h19C4] = 8'h00;
RAM[16'h19C5] = 8'h00;
RAM[16'h19C6] = 8'h00;
RAM[16'h19C7] = 8'h00;
RAM[16'h19C8] = 8'h00;
RAM[16'h19C9] = 8'h00;
RAM[16'h19CA] = 8'h00;
RAM[16'h19CB] = 8'h00;
RAM[16'h19CC] = 8'h00;
RAM[16'h19CD] = 8'h00;
RAM[16'h19CE] = 8'h00;
RAM[16'h19CF] = 8'h00;
RAM[16'h19D0] = 8'h00;
RAM[16'h19D1] = 8'h00;
RAM[16'h19D2] = 8'h00;
RAM[16'h19D3] = 8'h00;
RAM[16'h19D4] = 8'h00;
RAM[16'h19D5] = 8'h00;
RAM[16'h19D6] = 8'h00;
RAM[16'h19D7] = 8'h00;
RAM[16'h19D8] = 8'h00;
RAM[16'h19D9] = 8'h00;
RAM[16'h19DA] = 8'h00;
RAM[16'h19DB] = 8'h00;
RAM[16'h19DC] = 8'h00;
RAM[16'h19DD] = 8'h00;
RAM[16'h19DE] = 8'h00;
RAM[16'h19DF] = 8'h00;
RAM[16'h19E0] = 8'h00;
RAM[16'h19E1] = 8'h00;
RAM[16'h19E2] = 8'h00;
RAM[16'h19E3] = 8'h00;
RAM[16'h19E4] = 8'h00;
RAM[16'h19E5] = 8'h00;
RAM[16'h19E6] = 8'h00;
RAM[16'h19E7] = 8'h00;
RAM[16'h19E8] = 8'h00;
RAM[16'h19E9] = 8'h00;
RAM[16'h19EA] = 8'h00;
RAM[16'h19EB] = 8'h00;
RAM[16'h19EC] = 8'h00;
RAM[16'h19ED] = 8'h00;
RAM[16'h19EE] = 8'h00;
RAM[16'h19EF] = 8'h00;
RAM[16'h19F0] = 8'h00;
RAM[16'h19F1] = 8'h00;
RAM[16'h19F2] = 8'h00;
RAM[16'h19F3] = 8'h00;
RAM[16'h19F4] = 8'h00;
RAM[16'h19F5] = 8'h00;
RAM[16'h19F6] = 8'h00;
RAM[16'h19F7] = 8'h00;
RAM[16'h19F8] = 8'h00;
RAM[16'h19F9] = 8'h00;
RAM[16'h19FA] = 8'h00;
RAM[16'h19FB] = 8'h00;
RAM[16'h19FC] = 8'h00;
RAM[16'h19FD] = 8'h00;
RAM[16'h19FE] = 8'h00;
RAM[16'h19FF] = 8'h00;
RAM[16'h1A00] = 8'h00;
RAM[16'h1A01] = 8'h00;
RAM[16'h1A02] = 8'h00;
RAM[16'h1A03] = 8'h00;
RAM[16'h1A04] = 8'h00;
RAM[16'h1A05] = 8'h00;
RAM[16'h1A06] = 8'h00;
RAM[16'h1A07] = 8'h00;
RAM[16'h1A08] = 8'h00;
RAM[16'h1A09] = 8'h00;
RAM[16'h1A0A] = 8'h00;
RAM[16'h1A0B] = 8'h00;
RAM[16'h1A0C] = 8'h00;
RAM[16'h1A0D] = 8'h00;
RAM[16'h1A0E] = 8'h00;
RAM[16'h1A0F] = 8'h00;
RAM[16'h1A10] = 8'h00;
RAM[16'h1A11] = 8'h00;
RAM[16'h1A12] = 8'h00;
RAM[16'h1A13] = 8'h00;
RAM[16'h1A14] = 8'h00;
RAM[16'h1A15] = 8'h00;
RAM[16'h1A16] = 8'h00;
RAM[16'h1A17] = 8'h00;
RAM[16'h1A18] = 8'h00;
RAM[16'h1A19] = 8'h00;
RAM[16'h1A1A] = 8'h00;
RAM[16'h1A1B] = 8'h00;
RAM[16'h1A1C] = 8'h00;
RAM[16'h1A1D] = 8'h00;
RAM[16'h1A1E] = 8'h00;
RAM[16'h1A1F] = 8'h00;
RAM[16'h1A20] = 8'h00;
RAM[16'h1A21] = 8'h00;
RAM[16'h1A22] = 8'h00;
RAM[16'h1A23] = 8'h00;
RAM[16'h1A24] = 8'h00;
RAM[16'h1A25] = 8'h00;
RAM[16'h1A26] = 8'h00;
RAM[16'h1A27] = 8'h00;
RAM[16'h1A28] = 8'h00;
RAM[16'h1A29] = 8'h00;
RAM[16'h1A2A] = 8'h00;
RAM[16'h1A2B] = 8'h00;
RAM[16'h1A2C] = 8'h00;
RAM[16'h1A2D] = 8'h00;
RAM[16'h1A2E] = 8'h00;
RAM[16'h1A2F] = 8'h00;
RAM[16'h1A30] = 8'h00;
RAM[16'h1A31] = 8'h00;
RAM[16'h1A32] = 8'h00;
RAM[16'h1A33] = 8'h00;
RAM[16'h1A34] = 8'h00;
RAM[16'h1A35] = 8'h00;
RAM[16'h1A36] = 8'h00;
RAM[16'h1A37] = 8'h00;
RAM[16'h1A38] = 8'h00;
RAM[16'h1A39] = 8'h00;
RAM[16'h1A3A] = 8'h00;
RAM[16'h1A3B] = 8'h00;
RAM[16'h1A3C] = 8'h00;
RAM[16'h1A3D] = 8'h00;
RAM[16'h1A3E] = 8'h00;
RAM[16'h1A3F] = 8'h00;
RAM[16'h1A40] = 8'h00;
RAM[16'h1A41] = 8'h00;
RAM[16'h1A42] = 8'h00;
RAM[16'h1A43] = 8'h00;
RAM[16'h1A44] = 8'h00;
RAM[16'h1A45] = 8'h00;
RAM[16'h1A46] = 8'h00;
RAM[16'h1A47] = 8'h00;
RAM[16'h1A48] = 8'h00;
RAM[16'h1A49] = 8'h00;
RAM[16'h1A4A] = 8'h00;
RAM[16'h1A4B] = 8'h00;
RAM[16'h1A4C] = 8'h00;
RAM[16'h1A4D] = 8'h00;
RAM[16'h1A4E] = 8'h00;
RAM[16'h1A4F] = 8'h00;
RAM[16'h1A50] = 8'h00;
RAM[16'h1A51] = 8'h00;
RAM[16'h1A52] = 8'h00;
RAM[16'h1A53] = 8'h00;
RAM[16'h1A54] = 8'h00;
RAM[16'h1A55] = 8'h00;
RAM[16'h1A56] = 8'h00;
RAM[16'h1A57] = 8'h00;
RAM[16'h1A58] = 8'h00;
RAM[16'h1A59] = 8'h00;
RAM[16'h1A5A] = 8'h00;
RAM[16'h1A5B] = 8'h00;
RAM[16'h1A5C] = 8'h00;
RAM[16'h1A5D] = 8'h00;
RAM[16'h1A5E] = 8'h00;
RAM[16'h1A5F] = 8'h00;
RAM[16'h1A60] = 8'h00;
RAM[16'h1A61] = 8'h00;
RAM[16'h1A62] = 8'h00;
RAM[16'h1A63] = 8'h00;
RAM[16'h1A64] = 8'h00;
RAM[16'h1A65] = 8'h00;
RAM[16'h1A66] = 8'h00;
RAM[16'h1A67] = 8'h00;
RAM[16'h1A68] = 8'h00;
RAM[16'h1A69] = 8'h00;
RAM[16'h1A6A] = 8'h00;
RAM[16'h1A6B] = 8'h00;
RAM[16'h1A6C] = 8'h00;
RAM[16'h1A6D] = 8'h00;
RAM[16'h1A6E] = 8'h00;
RAM[16'h1A6F] = 8'h00;
RAM[16'h1A70] = 8'h00;
RAM[16'h1A71] = 8'h00;
RAM[16'h1A72] = 8'h00;
RAM[16'h1A73] = 8'h00;
RAM[16'h1A74] = 8'h00;
RAM[16'h1A75] = 8'h00;
RAM[16'h1A76] = 8'h00;
RAM[16'h1A77] = 8'h00;
RAM[16'h1A78] = 8'h00;
RAM[16'h1A79] = 8'h00;
RAM[16'h1A7A] = 8'h00;
RAM[16'h1A7B] = 8'h00;
RAM[16'h1A7C] = 8'h00;
RAM[16'h1A7D] = 8'h00;
RAM[16'h1A7E] = 8'h00;
RAM[16'h1A7F] = 8'h00;
RAM[16'h1A80] = 8'h00;
RAM[16'h1A81] = 8'h00;
RAM[16'h1A82] = 8'h00;
RAM[16'h1A83] = 8'h00;
RAM[16'h1A84] = 8'h00;
RAM[16'h1A85] = 8'h00;
RAM[16'h1A86] = 8'h00;
RAM[16'h1A87] = 8'h00;
RAM[16'h1A88] = 8'h00;
RAM[16'h1A89] = 8'h00;
RAM[16'h1A8A] = 8'h00;
RAM[16'h1A8B] = 8'h00;
RAM[16'h1A8C] = 8'h00;
RAM[16'h1A8D] = 8'h00;
RAM[16'h1A8E] = 8'h00;
RAM[16'h1A8F] = 8'h00;
RAM[16'h1A90] = 8'h00;
RAM[16'h1A91] = 8'h00;
RAM[16'h1A92] = 8'h00;
RAM[16'h1A93] = 8'h00;
RAM[16'h1A94] = 8'h00;
RAM[16'h1A95] = 8'h00;
RAM[16'h1A96] = 8'h00;
RAM[16'h1A97] = 8'h00;
RAM[16'h1A98] = 8'h00;
RAM[16'h1A99] = 8'h00;
RAM[16'h1A9A] = 8'h00;
RAM[16'h1A9B] = 8'h00;
RAM[16'h1A9C] = 8'h00;
RAM[16'h1A9D] = 8'h00;
RAM[16'h1A9E] = 8'h00;
RAM[16'h1A9F] = 8'h00;
RAM[16'h1AA0] = 8'h00;
RAM[16'h1AA1] = 8'h00;
RAM[16'h1AA2] = 8'h00;
RAM[16'h1AA3] = 8'h00;
RAM[16'h1AA4] = 8'h00;
RAM[16'h1AA5] = 8'h00;
RAM[16'h1AA6] = 8'h00;
RAM[16'h1AA7] = 8'h00;
RAM[16'h1AA8] = 8'h00;
RAM[16'h1AA9] = 8'h00;
RAM[16'h1AAA] = 8'h00;
RAM[16'h1AAB] = 8'h00;
RAM[16'h1AAC] = 8'h00;
RAM[16'h1AAD] = 8'h00;
RAM[16'h1AAE] = 8'h00;
RAM[16'h1AAF] = 8'h00;
RAM[16'h1AB0] = 8'h00;
RAM[16'h1AB1] = 8'h00;
RAM[16'h1AB2] = 8'h00;
RAM[16'h1AB3] = 8'h00;
RAM[16'h1AB4] = 8'h00;
RAM[16'h1AB5] = 8'h00;
RAM[16'h1AB6] = 8'h00;
RAM[16'h1AB7] = 8'h00;
RAM[16'h1AB8] = 8'h00;
RAM[16'h1AB9] = 8'h00;
RAM[16'h1ABA] = 8'h00;
RAM[16'h1ABB] = 8'h00;
RAM[16'h1ABC] = 8'h00;
RAM[16'h1ABD] = 8'h00;
RAM[16'h1ABE] = 8'h00;
RAM[16'h1ABF] = 8'h00;
RAM[16'h1AC0] = 8'h00;
RAM[16'h1AC1] = 8'h00;
RAM[16'h1AC2] = 8'h00;
RAM[16'h1AC3] = 8'h00;
RAM[16'h1AC4] = 8'h00;
RAM[16'h1AC5] = 8'h00;
RAM[16'h1AC6] = 8'h00;
RAM[16'h1AC7] = 8'h00;
RAM[16'h1AC8] = 8'h00;
RAM[16'h1AC9] = 8'h00;
RAM[16'h1ACA] = 8'h00;
RAM[16'h1ACB] = 8'h00;
RAM[16'h1ACC] = 8'h00;
RAM[16'h1ACD] = 8'h00;
RAM[16'h1ACE] = 8'h00;
RAM[16'h1ACF] = 8'h00;
RAM[16'h1AD0] = 8'h00;
RAM[16'h1AD1] = 8'h00;
RAM[16'h1AD2] = 8'h00;
RAM[16'h1AD3] = 8'h00;
RAM[16'h1AD4] = 8'h00;
RAM[16'h1AD5] = 8'h00;
RAM[16'h1AD6] = 8'h00;
RAM[16'h1AD7] = 8'h00;
RAM[16'h1AD8] = 8'h00;
RAM[16'h1AD9] = 8'h00;
RAM[16'h1ADA] = 8'h00;
RAM[16'h1ADB] = 8'h00;
RAM[16'h1ADC] = 8'h00;
RAM[16'h1ADD] = 8'h00;
RAM[16'h1ADE] = 8'h00;
RAM[16'h1ADF] = 8'h00;
RAM[16'h1AE0] = 8'h00;
RAM[16'h1AE1] = 8'h00;
RAM[16'h1AE2] = 8'h00;
RAM[16'h1AE3] = 8'h00;
RAM[16'h1AE4] = 8'h00;
RAM[16'h1AE5] = 8'h00;
RAM[16'h1AE6] = 8'h00;
RAM[16'h1AE7] = 8'h00;
RAM[16'h1AE8] = 8'h00;
RAM[16'h1AE9] = 8'h00;
RAM[16'h1AEA] = 8'h00;
RAM[16'h1AEB] = 8'h00;
RAM[16'h1AEC] = 8'h00;
RAM[16'h1AED] = 8'h00;
RAM[16'h1AEE] = 8'h00;
RAM[16'h1AEF] = 8'h00;
RAM[16'h1AF0] = 8'h00;
RAM[16'h1AF1] = 8'h00;
RAM[16'h1AF2] = 8'h00;
RAM[16'h1AF3] = 8'h00;
RAM[16'h1AF4] = 8'h00;
RAM[16'h1AF5] = 8'h00;
RAM[16'h1AF6] = 8'h00;
RAM[16'h1AF7] = 8'h00;
RAM[16'h1AF8] = 8'h00;
RAM[16'h1AF9] = 8'h00;
RAM[16'h1AFA] = 8'h00;
RAM[16'h1AFB] = 8'h00;
RAM[16'h1AFC] = 8'h00;
RAM[16'h1AFD] = 8'h00;
RAM[16'h1AFE] = 8'h00;
RAM[16'h1AFF] = 8'h00;
RAM[16'h1B00] = 8'h00;
RAM[16'h1B01] = 8'h00;
RAM[16'h1B02] = 8'h00;
RAM[16'h1B03] = 8'h00;
RAM[16'h1B04] = 8'h00;
RAM[16'h1B05] = 8'h00;
RAM[16'h1B06] = 8'h00;
RAM[16'h1B07] = 8'h00;
RAM[16'h1B08] = 8'h00;
RAM[16'h1B09] = 8'h00;
RAM[16'h1B0A] = 8'h00;
RAM[16'h1B0B] = 8'h00;
RAM[16'h1B0C] = 8'h00;
RAM[16'h1B0D] = 8'h00;
RAM[16'h1B0E] = 8'h00;
RAM[16'h1B0F] = 8'h00;
RAM[16'h1B10] = 8'h00;
RAM[16'h1B11] = 8'h00;
RAM[16'h1B12] = 8'h00;
RAM[16'h1B13] = 8'h00;
RAM[16'h1B14] = 8'h00;
RAM[16'h1B15] = 8'h00;
RAM[16'h1B16] = 8'h00;
RAM[16'h1B17] = 8'h00;
RAM[16'h1B18] = 8'h00;
RAM[16'h1B19] = 8'h00;
RAM[16'h1B1A] = 8'h00;
RAM[16'h1B1B] = 8'h00;
RAM[16'h1B1C] = 8'h00;
RAM[16'h1B1D] = 8'h00;
RAM[16'h1B1E] = 8'h00;
RAM[16'h1B1F] = 8'h00;
RAM[16'h1B20] = 8'h00;
RAM[16'h1B21] = 8'h00;
RAM[16'h1B22] = 8'h00;
RAM[16'h1B23] = 8'h00;
RAM[16'h1B24] = 8'h00;
RAM[16'h1B25] = 8'h00;
RAM[16'h1B26] = 8'h00;
RAM[16'h1B27] = 8'h00;
RAM[16'h1B28] = 8'h00;
RAM[16'h1B29] = 8'h00;
RAM[16'h1B2A] = 8'h00;
RAM[16'h1B2B] = 8'h00;
RAM[16'h1B2C] = 8'h00;
RAM[16'h1B2D] = 8'h00;
RAM[16'h1B2E] = 8'h00;
RAM[16'h1B2F] = 8'h00;
RAM[16'h1B30] = 8'h00;
RAM[16'h1B31] = 8'h00;
RAM[16'h1B32] = 8'h00;
RAM[16'h1B33] = 8'h00;
RAM[16'h1B34] = 8'h00;
RAM[16'h1B35] = 8'h00;
RAM[16'h1B36] = 8'h00;
RAM[16'h1B37] = 8'h00;
RAM[16'h1B38] = 8'h00;
RAM[16'h1B39] = 8'h00;
RAM[16'h1B3A] = 8'h00;
RAM[16'h1B3B] = 8'h00;
RAM[16'h1B3C] = 8'h00;
RAM[16'h1B3D] = 8'h00;
RAM[16'h1B3E] = 8'h00;
RAM[16'h1B3F] = 8'h00;
RAM[16'h1B40] = 8'h00;
RAM[16'h1B41] = 8'h00;
RAM[16'h1B42] = 8'h00;
RAM[16'h1B43] = 8'h00;
RAM[16'h1B44] = 8'h00;
RAM[16'h1B45] = 8'h00;
RAM[16'h1B46] = 8'h00;
RAM[16'h1B47] = 8'h00;
RAM[16'h1B48] = 8'h00;
RAM[16'h1B49] = 8'h00;
RAM[16'h1B4A] = 8'h00;
RAM[16'h1B4B] = 8'h00;
RAM[16'h1B4C] = 8'h00;
RAM[16'h1B4D] = 8'h00;
RAM[16'h1B4E] = 8'h00;
RAM[16'h1B4F] = 8'h00;
RAM[16'h1B50] = 8'h00;
RAM[16'h1B51] = 8'h00;
RAM[16'h1B52] = 8'h00;
RAM[16'h1B53] = 8'h00;
RAM[16'h1B54] = 8'h00;
RAM[16'h1B55] = 8'h00;
RAM[16'h1B56] = 8'h00;
RAM[16'h1B57] = 8'h00;
RAM[16'h1B58] = 8'h00;
RAM[16'h1B59] = 8'h00;
RAM[16'h1B5A] = 8'h00;
RAM[16'h1B5B] = 8'h00;
RAM[16'h1B5C] = 8'h00;
RAM[16'h1B5D] = 8'h00;
RAM[16'h1B5E] = 8'h00;
RAM[16'h1B5F] = 8'h00;
RAM[16'h1B60] = 8'h00;
RAM[16'h1B61] = 8'h00;
RAM[16'h1B62] = 8'h00;
RAM[16'h1B63] = 8'h00;
RAM[16'h1B64] = 8'h00;
RAM[16'h1B65] = 8'h00;
RAM[16'h1B66] = 8'h00;
RAM[16'h1B67] = 8'h00;
RAM[16'h1B68] = 8'h00;
RAM[16'h1B69] = 8'h00;
RAM[16'h1B6A] = 8'h00;
RAM[16'h1B6B] = 8'h00;
RAM[16'h1B6C] = 8'h00;
RAM[16'h1B6D] = 8'h00;
RAM[16'h1B6E] = 8'h00;
RAM[16'h1B6F] = 8'h00;
RAM[16'h1B70] = 8'h00;
RAM[16'h1B71] = 8'h00;
RAM[16'h1B72] = 8'h00;
RAM[16'h1B73] = 8'h00;
RAM[16'h1B74] = 8'h00;
RAM[16'h1B75] = 8'h00;
RAM[16'h1B76] = 8'h00;
RAM[16'h1B77] = 8'h00;
RAM[16'h1B78] = 8'h00;
RAM[16'h1B79] = 8'h00;
RAM[16'h1B7A] = 8'h00;
RAM[16'h1B7B] = 8'h00;
RAM[16'h1B7C] = 8'h00;
RAM[16'h1B7D] = 8'h00;
RAM[16'h1B7E] = 8'h00;
RAM[16'h1B7F] = 8'h00;
RAM[16'h1B80] = 8'h00;
RAM[16'h1B81] = 8'h00;
RAM[16'h1B82] = 8'h00;
RAM[16'h1B83] = 8'h00;
RAM[16'h1B84] = 8'h00;
RAM[16'h1B85] = 8'h00;
RAM[16'h1B86] = 8'h00;
RAM[16'h1B87] = 8'h00;
RAM[16'h1B88] = 8'h00;
RAM[16'h1B89] = 8'h00;
RAM[16'h1B8A] = 8'h00;
RAM[16'h1B8B] = 8'h00;
RAM[16'h1B8C] = 8'h00;
RAM[16'h1B8D] = 8'h00;
RAM[16'h1B8E] = 8'h00;
RAM[16'h1B8F] = 8'h00;
RAM[16'h1B90] = 8'h00;
RAM[16'h1B91] = 8'h00;
RAM[16'h1B92] = 8'h00;
RAM[16'h1B93] = 8'h00;
RAM[16'h1B94] = 8'h00;
RAM[16'h1B95] = 8'h00;
RAM[16'h1B96] = 8'h00;
RAM[16'h1B97] = 8'h00;
RAM[16'h1B98] = 8'h00;
RAM[16'h1B99] = 8'h00;
RAM[16'h1B9A] = 8'h00;
RAM[16'h1B9B] = 8'h00;
RAM[16'h1B9C] = 8'h00;
RAM[16'h1B9D] = 8'h00;
RAM[16'h1B9E] = 8'h00;
RAM[16'h1B9F] = 8'h00;
RAM[16'h1BA0] = 8'h00;
RAM[16'h1BA1] = 8'h00;
RAM[16'h1BA2] = 8'h00;
RAM[16'h1BA3] = 8'h00;
RAM[16'h1BA4] = 8'h00;
RAM[16'h1BA5] = 8'h00;
RAM[16'h1BA6] = 8'h00;
RAM[16'h1BA7] = 8'h00;
RAM[16'h1BA8] = 8'h00;
RAM[16'h1BA9] = 8'h00;
RAM[16'h1BAA] = 8'h00;
RAM[16'h1BAB] = 8'h00;
RAM[16'h1BAC] = 8'h00;
RAM[16'h1BAD] = 8'h00;
RAM[16'h1BAE] = 8'h00;
RAM[16'h1BAF] = 8'h00;
RAM[16'h1BB0] = 8'h00;
RAM[16'h1BB1] = 8'h00;
RAM[16'h1BB2] = 8'h00;
RAM[16'h1BB3] = 8'h00;
RAM[16'h1BB4] = 8'h00;
RAM[16'h1BB5] = 8'h00;
RAM[16'h1BB6] = 8'h00;
RAM[16'h1BB7] = 8'h00;
RAM[16'h1BB8] = 8'h00;
RAM[16'h1BB9] = 8'h00;
RAM[16'h1BBA] = 8'h00;
RAM[16'h1BBB] = 8'h00;
RAM[16'h1BBC] = 8'h00;
RAM[16'h1BBD] = 8'h00;
RAM[16'h1BBE] = 8'h00;
RAM[16'h1BBF] = 8'h00;
RAM[16'h1BC0] = 8'h00;
RAM[16'h1BC1] = 8'h00;
RAM[16'h1BC2] = 8'h00;
RAM[16'h1BC3] = 8'h00;
RAM[16'h1BC4] = 8'h00;
RAM[16'h1BC5] = 8'h00;
RAM[16'h1BC6] = 8'h00;
RAM[16'h1BC7] = 8'h00;
RAM[16'h1BC8] = 8'h00;
RAM[16'h1BC9] = 8'h00;
RAM[16'h1BCA] = 8'h00;
RAM[16'h1BCB] = 8'h00;
RAM[16'h1BCC] = 8'h00;
RAM[16'h1BCD] = 8'h00;
RAM[16'h1BCE] = 8'h00;
RAM[16'h1BCF] = 8'h00;
RAM[16'h1BD0] = 8'h00;
RAM[16'h1BD1] = 8'h00;
RAM[16'h1BD2] = 8'h00;
RAM[16'h1BD3] = 8'h00;
RAM[16'h1BD4] = 8'h00;
RAM[16'h1BD5] = 8'h00;
RAM[16'h1BD6] = 8'h00;
RAM[16'h1BD7] = 8'h00;
RAM[16'h1BD8] = 8'h00;
RAM[16'h1BD9] = 8'h00;
RAM[16'h1BDA] = 8'h00;
RAM[16'h1BDB] = 8'h00;
RAM[16'h1BDC] = 8'h00;
RAM[16'h1BDD] = 8'h00;
RAM[16'h1BDE] = 8'h00;
RAM[16'h1BDF] = 8'h00;
RAM[16'h1BE0] = 8'h00;
RAM[16'h1BE1] = 8'h00;
RAM[16'h1BE2] = 8'h00;
RAM[16'h1BE3] = 8'h00;
RAM[16'h1BE4] = 8'h00;
RAM[16'h1BE5] = 8'h00;
RAM[16'h1BE6] = 8'h00;
RAM[16'h1BE7] = 8'h00;
RAM[16'h1BE8] = 8'h00;
RAM[16'h1BE9] = 8'h00;
RAM[16'h1BEA] = 8'h00;
RAM[16'h1BEB] = 8'h00;
RAM[16'h1BEC] = 8'h00;
RAM[16'h1BED] = 8'h00;
RAM[16'h1BEE] = 8'h00;
RAM[16'h1BEF] = 8'h00;
RAM[16'h1BF0] = 8'h00;
RAM[16'h1BF1] = 8'h00;
RAM[16'h1BF2] = 8'h00;
RAM[16'h1BF3] = 8'h00;
RAM[16'h1BF4] = 8'h00;
RAM[16'h1BF5] = 8'h00;
RAM[16'h1BF6] = 8'h00;
RAM[16'h1BF7] = 8'h00;
RAM[16'h1BF8] = 8'h00;
RAM[16'h1BF9] = 8'h00;
RAM[16'h1BFA] = 8'h00;
RAM[16'h1BFB] = 8'h00;
RAM[16'h1BFC] = 8'h00;
RAM[16'h1BFD] = 8'h00;
RAM[16'h1BFE] = 8'h00;
RAM[16'h1BFF] = 8'h00;
RAM[16'h1C00] = 8'h00;
RAM[16'h1C01] = 8'h00;
RAM[16'h1C02] = 8'h00;
RAM[16'h1C03] = 8'h00;
RAM[16'h1C04] = 8'h00;
RAM[16'h1C05] = 8'h00;
RAM[16'h1C06] = 8'h00;
RAM[16'h1C07] = 8'h00;
RAM[16'h1C08] = 8'h00;
RAM[16'h1C09] = 8'h00;
RAM[16'h1C0A] = 8'h00;
RAM[16'h1C0B] = 8'h00;
RAM[16'h1C0C] = 8'h00;
RAM[16'h1C0D] = 8'h00;
RAM[16'h1C0E] = 8'h00;
RAM[16'h1C0F] = 8'h00;
RAM[16'h1C10] = 8'h00;
RAM[16'h1C11] = 8'h00;
RAM[16'h1C12] = 8'h00;
RAM[16'h1C13] = 8'h00;
RAM[16'h1C14] = 8'h00;
RAM[16'h1C15] = 8'h00;
RAM[16'h1C16] = 8'h00;
RAM[16'h1C17] = 8'h00;
RAM[16'h1C18] = 8'h00;
RAM[16'h1C19] = 8'h00;
RAM[16'h1C1A] = 8'h00;
RAM[16'h1C1B] = 8'h00;
RAM[16'h1C1C] = 8'h00;
RAM[16'h1C1D] = 8'h00;
RAM[16'h1C1E] = 8'h00;
RAM[16'h1C1F] = 8'h00;
RAM[16'h1C20] = 8'h00;
RAM[16'h1C21] = 8'h00;
RAM[16'h1C22] = 8'h00;
RAM[16'h1C23] = 8'h00;
RAM[16'h1C24] = 8'h00;
RAM[16'h1C25] = 8'h00;
RAM[16'h1C26] = 8'h00;
RAM[16'h1C27] = 8'h00;
RAM[16'h1C28] = 8'h00;
RAM[16'h1C29] = 8'h00;
RAM[16'h1C2A] = 8'h00;
RAM[16'h1C2B] = 8'h00;
RAM[16'h1C2C] = 8'h00;
RAM[16'h1C2D] = 8'h00;
RAM[16'h1C2E] = 8'h00;
RAM[16'h1C2F] = 8'h00;
RAM[16'h1C30] = 8'h00;
RAM[16'h1C31] = 8'h00;
RAM[16'h1C32] = 8'h00;
RAM[16'h1C33] = 8'h00;
RAM[16'h1C34] = 8'h00;
RAM[16'h1C35] = 8'h00;
RAM[16'h1C36] = 8'h00;
RAM[16'h1C37] = 8'h00;
RAM[16'h1C38] = 8'h00;
RAM[16'h1C39] = 8'h00;
RAM[16'h1C3A] = 8'h00;
RAM[16'h1C3B] = 8'h00;
RAM[16'h1C3C] = 8'h00;
RAM[16'h1C3D] = 8'h00;
RAM[16'h1C3E] = 8'h00;
RAM[16'h1C3F] = 8'h00;
RAM[16'h1C40] = 8'h00;
RAM[16'h1C41] = 8'h00;
RAM[16'h1C42] = 8'h00;
RAM[16'h1C43] = 8'h00;
RAM[16'h1C44] = 8'h00;
RAM[16'h1C45] = 8'h00;
RAM[16'h1C46] = 8'h00;
RAM[16'h1C47] = 8'h00;
RAM[16'h1C48] = 8'h00;
RAM[16'h1C49] = 8'h00;
RAM[16'h1C4A] = 8'h00;
RAM[16'h1C4B] = 8'h00;
RAM[16'h1C4C] = 8'h00;
RAM[16'h1C4D] = 8'h00;
RAM[16'h1C4E] = 8'h00;
RAM[16'h1C4F] = 8'h00;
RAM[16'h1C50] = 8'h00;
RAM[16'h1C51] = 8'h00;
RAM[16'h1C52] = 8'h00;
RAM[16'h1C53] = 8'h00;
RAM[16'h1C54] = 8'h00;
RAM[16'h1C55] = 8'h00;
RAM[16'h1C56] = 8'h00;
RAM[16'h1C57] = 8'h00;
RAM[16'h1C58] = 8'h00;
RAM[16'h1C59] = 8'h00;
RAM[16'h1C5A] = 8'h00;
RAM[16'h1C5B] = 8'h00;
RAM[16'h1C5C] = 8'h00;
RAM[16'h1C5D] = 8'h00;
RAM[16'h1C5E] = 8'h00;
RAM[16'h1C5F] = 8'h00;
RAM[16'h1C60] = 8'h00;
RAM[16'h1C61] = 8'h00;
RAM[16'h1C62] = 8'h00;
RAM[16'h1C63] = 8'h00;
RAM[16'h1C64] = 8'h00;
RAM[16'h1C65] = 8'h00;
RAM[16'h1C66] = 8'h00;
RAM[16'h1C67] = 8'h00;
RAM[16'h1C68] = 8'h00;
RAM[16'h1C69] = 8'h00;
RAM[16'h1C6A] = 8'h00;
RAM[16'h1C6B] = 8'h00;
RAM[16'h1C6C] = 8'h00;
RAM[16'h1C6D] = 8'h00;
RAM[16'h1C6E] = 8'h00;
RAM[16'h1C6F] = 8'h00;
RAM[16'h1C70] = 8'h00;
RAM[16'h1C71] = 8'h00;
RAM[16'h1C72] = 8'h00;
RAM[16'h1C73] = 8'h00;
RAM[16'h1C74] = 8'h00;
RAM[16'h1C75] = 8'h00;
RAM[16'h1C76] = 8'h00;
RAM[16'h1C77] = 8'h00;
RAM[16'h1C78] = 8'h00;
RAM[16'h1C79] = 8'h00;
RAM[16'h1C7A] = 8'h00;
RAM[16'h1C7B] = 8'h00;
RAM[16'h1C7C] = 8'h00;
RAM[16'h1C7D] = 8'h00;
RAM[16'h1C7E] = 8'h00;
RAM[16'h1C7F] = 8'h00;
RAM[16'h1C80] = 8'h00;
RAM[16'h1C81] = 8'h00;
RAM[16'h1C82] = 8'h00;
RAM[16'h1C83] = 8'h00;
RAM[16'h1C84] = 8'h00;
RAM[16'h1C85] = 8'h00;
RAM[16'h1C86] = 8'h00;
RAM[16'h1C87] = 8'h00;
RAM[16'h1C88] = 8'h00;
RAM[16'h1C89] = 8'h00;
RAM[16'h1C8A] = 8'h00;
RAM[16'h1C8B] = 8'h00;
RAM[16'h1C8C] = 8'h00;
RAM[16'h1C8D] = 8'h00;
RAM[16'h1C8E] = 8'h00;
RAM[16'h1C8F] = 8'h00;
RAM[16'h1C90] = 8'h00;
RAM[16'h1C91] = 8'h00;
RAM[16'h1C92] = 8'h00;
RAM[16'h1C93] = 8'h00;
RAM[16'h1C94] = 8'h00;
RAM[16'h1C95] = 8'h00;
RAM[16'h1C96] = 8'h00;
RAM[16'h1C97] = 8'h00;
RAM[16'h1C98] = 8'h00;
RAM[16'h1C99] = 8'h00;
RAM[16'h1C9A] = 8'h00;
RAM[16'h1C9B] = 8'h00;
RAM[16'h1C9C] = 8'h00;
RAM[16'h1C9D] = 8'h00;
RAM[16'h1C9E] = 8'h00;
RAM[16'h1C9F] = 8'h00;
RAM[16'h1CA0] = 8'h00;
RAM[16'h1CA1] = 8'h00;
RAM[16'h1CA2] = 8'h00;
RAM[16'h1CA3] = 8'h00;
RAM[16'h1CA4] = 8'h00;
RAM[16'h1CA5] = 8'h00;
RAM[16'h1CA6] = 8'h00;
RAM[16'h1CA7] = 8'h00;
RAM[16'h1CA8] = 8'h00;
RAM[16'h1CA9] = 8'h00;
RAM[16'h1CAA] = 8'h00;
RAM[16'h1CAB] = 8'h00;
RAM[16'h1CAC] = 8'h00;
RAM[16'h1CAD] = 8'h00;
RAM[16'h1CAE] = 8'h00;
RAM[16'h1CAF] = 8'h00;
RAM[16'h1CB0] = 8'h00;
RAM[16'h1CB1] = 8'h00;
RAM[16'h1CB2] = 8'h00;
RAM[16'h1CB3] = 8'h00;
RAM[16'h1CB4] = 8'h00;
RAM[16'h1CB5] = 8'h00;
RAM[16'h1CB6] = 8'h00;
RAM[16'h1CB7] = 8'h00;
RAM[16'h1CB8] = 8'h00;
RAM[16'h1CB9] = 8'h00;
RAM[16'h1CBA] = 8'h00;
RAM[16'h1CBB] = 8'h00;
RAM[16'h1CBC] = 8'h00;
RAM[16'h1CBD] = 8'h00;
RAM[16'h1CBE] = 8'h00;
RAM[16'h1CBF] = 8'h00;
RAM[16'h1CC0] = 8'h00;
RAM[16'h1CC1] = 8'h00;
RAM[16'h1CC2] = 8'h00;
RAM[16'h1CC3] = 8'h00;
RAM[16'h1CC4] = 8'h00;
RAM[16'h1CC5] = 8'h00;
RAM[16'h1CC6] = 8'h00;
RAM[16'h1CC7] = 8'h00;
RAM[16'h1CC8] = 8'h00;
RAM[16'h1CC9] = 8'h00;
RAM[16'h1CCA] = 8'h00;
RAM[16'h1CCB] = 8'h00;
RAM[16'h1CCC] = 8'h00;
RAM[16'h1CCD] = 8'h00;
RAM[16'h1CCE] = 8'h00;
RAM[16'h1CCF] = 8'h00;
RAM[16'h1CD0] = 8'h00;
RAM[16'h1CD1] = 8'h00;
RAM[16'h1CD2] = 8'h00;
RAM[16'h1CD3] = 8'h00;
RAM[16'h1CD4] = 8'h00;
RAM[16'h1CD5] = 8'h00;
RAM[16'h1CD6] = 8'h00;
RAM[16'h1CD7] = 8'h00;
RAM[16'h1CD8] = 8'h00;
RAM[16'h1CD9] = 8'h00;
RAM[16'h1CDA] = 8'h00;
RAM[16'h1CDB] = 8'h00;
RAM[16'h1CDC] = 8'h00;
RAM[16'h1CDD] = 8'h00;
RAM[16'h1CDE] = 8'h00;
RAM[16'h1CDF] = 8'h00;
RAM[16'h1CE0] = 8'h00;
RAM[16'h1CE1] = 8'h00;
RAM[16'h1CE2] = 8'h00;
RAM[16'h1CE3] = 8'h00;
RAM[16'h1CE4] = 8'h00;
RAM[16'h1CE5] = 8'h00;
RAM[16'h1CE6] = 8'h00;
RAM[16'h1CE7] = 8'h00;
RAM[16'h1CE8] = 8'h00;
RAM[16'h1CE9] = 8'h00;
RAM[16'h1CEA] = 8'h00;
RAM[16'h1CEB] = 8'h00;
RAM[16'h1CEC] = 8'h00;
RAM[16'h1CED] = 8'h00;
RAM[16'h1CEE] = 8'h00;
RAM[16'h1CEF] = 8'h00;
RAM[16'h1CF0] = 8'h00;
RAM[16'h1CF1] = 8'h00;
RAM[16'h1CF2] = 8'h00;
RAM[16'h1CF3] = 8'h00;
RAM[16'h1CF4] = 8'h00;
RAM[16'h1CF5] = 8'h00;
RAM[16'h1CF6] = 8'h00;
RAM[16'h1CF7] = 8'h00;
RAM[16'h1CF8] = 8'h00;
RAM[16'h1CF9] = 8'h00;
RAM[16'h1CFA] = 8'h00;
RAM[16'h1CFB] = 8'h00;
RAM[16'h1CFC] = 8'h00;
RAM[16'h1CFD] = 8'h00;
RAM[16'h1CFE] = 8'h00;
RAM[16'h1CFF] = 8'h00;
RAM[16'h1D00] = 8'h00;
RAM[16'h1D01] = 8'h00;
RAM[16'h1D02] = 8'h00;
RAM[16'h1D03] = 8'h00;
RAM[16'h1D04] = 8'h00;
RAM[16'h1D05] = 8'h00;
RAM[16'h1D06] = 8'h00;
RAM[16'h1D07] = 8'h00;
RAM[16'h1D08] = 8'h00;
RAM[16'h1D09] = 8'h00;
RAM[16'h1D0A] = 8'h00;
RAM[16'h1D0B] = 8'h00;
RAM[16'h1D0C] = 8'h00;
RAM[16'h1D0D] = 8'h00;
RAM[16'h1D0E] = 8'h00;
RAM[16'h1D0F] = 8'h00;
RAM[16'h1D10] = 8'h00;
RAM[16'h1D11] = 8'h00;
RAM[16'h1D12] = 8'h00;
RAM[16'h1D13] = 8'h00;
RAM[16'h1D14] = 8'h00;
RAM[16'h1D15] = 8'h00;
RAM[16'h1D16] = 8'h00;
RAM[16'h1D17] = 8'h00;
RAM[16'h1D18] = 8'h00;
RAM[16'h1D19] = 8'h00;
RAM[16'h1D1A] = 8'h00;
RAM[16'h1D1B] = 8'h00;
RAM[16'h1D1C] = 8'h00;
RAM[16'h1D1D] = 8'h00;
RAM[16'h1D1E] = 8'h00;
RAM[16'h1D1F] = 8'h00;
RAM[16'h1D20] = 8'h00;
RAM[16'h1D21] = 8'h00;
RAM[16'h1D22] = 8'h00;
RAM[16'h1D23] = 8'h00;
RAM[16'h1D24] = 8'h00;
RAM[16'h1D25] = 8'h00;
RAM[16'h1D26] = 8'h00;
RAM[16'h1D27] = 8'h00;
RAM[16'h1D28] = 8'h00;
RAM[16'h1D29] = 8'h00;
RAM[16'h1D2A] = 8'h00;
RAM[16'h1D2B] = 8'h00;
RAM[16'h1D2C] = 8'h00;
RAM[16'h1D2D] = 8'h00;
RAM[16'h1D2E] = 8'h00;
RAM[16'h1D2F] = 8'h00;
RAM[16'h1D30] = 8'h00;
RAM[16'h1D31] = 8'h00;
RAM[16'h1D32] = 8'h00;
RAM[16'h1D33] = 8'h00;
RAM[16'h1D34] = 8'h00;
RAM[16'h1D35] = 8'h00;
RAM[16'h1D36] = 8'h00;
RAM[16'h1D37] = 8'h00;
RAM[16'h1D38] = 8'h00;
RAM[16'h1D39] = 8'h00;
RAM[16'h1D3A] = 8'h00;
RAM[16'h1D3B] = 8'h00;
RAM[16'h1D3C] = 8'h00;
RAM[16'h1D3D] = 8'h00;
RAM[16'h1D3E] = 8'h00;
RAM[16'h1D3F] = 8'h00;
RAM[16'h1D40] = 8'h00;
RAM[16'h1D41] = 8'h00;
RAM[16'h1D42] = 8'h00;
RAM[16'h1D43] = 8'h00;
RAM[16'h1D44] = 8'h00;
RAM[16'h1D45] = 8'h00;
RAM[16'h1D46] = 8'h00;
RAM[16'h1D47] = 8'h00;
RAM[16'h1D48] = 8'h00;
RAM[16'h1D49] = 8'h00;
RAM[16'h1D4A] = 8'h00;
RAM[16'h1D4B] = 8'h00;
RAM[16'h1D4C] = 8'h00;
RAM[16'h1D4D] = 8'h00;
RAM[16'h1D4E] = 8'h00;
RAM[16'h1D4F] = 8'h00;
RAM[16'h1D50] = 8'h00;
RAM[16'h1D51] = 8'h00;
RAM[16'h1D52] = 8'h00;
RAM[16'h1D53] = 8'h00;
RAM[16'h1D54] = 8'h00;
RAM[16'h1D55] = 8'h00;
RAM[16'h1D56] = 8'h00;
RAM[16'h1D57] = 8'h00;
RAM[16'h1D58] = 8'h00;
RAM[16'h1D59] = 8'h00;
RAM[16'h1D5A] = 8'h00;
RAM[16'h1D5B] = 8'h00;
RAM[16'h1D5C] = 8'h00;
RAM[16'h1D5D] = 8'h00;
RAM[16'h1D5E] = 8'h00;
RAM[16'h1D5F] = 8'h00;
RAM[16'h1D60] = 8'h00;
RAM[16'h1D61] = 8'h00;
RAM[16'h1D62] = 8'h00;
RAM[16'h1D63] = 8'h00;
RAM[16'h1D64] = 8'h00;
RAM[16'h1D65] = 8'h00;
RAM[16'h1D66] = 8'h00;
RAM[16'h1D67] = 8'h00;
RAM[16'h1D68] = 8'h00;
RAM[16'h1D69] = 8'h00;
RAM[16'h1D6A] = 8'h00;
RAM[16'h1D6B] = 8'h00;
RAM[16'h1D6C] = 8'h00;
RAM[16'h1D6D] = 8'h00;
RAM[16'h1D6E] = 8'h00;
RAM[16'h1D6F] = 8'h00;
RAM[16'h1D70] = 8'h00;
RAM[16'h1D71] = 8'h00;
RAM[16'h1D72] = 8'h00;
RAM[16'h1D73] = 8'h00;
RAM[16'h1D74] = 8'h00;
RAM[16'h1D75] = 8'h00;
RAM[16'h1D76] = 8'h00;
RAM[16'h1D77] = 8'h00;
RAM[16'h1D78] = 8'h00;
RAM[16'h1D79] = 8'h00;
RAM[16'h1D7A] = 8'h00;
RAM[16'h1D7B] = 8'h00;
RAM[16'h1D7C] = 8'h00;
RAM[16'h1D7D] = 8'h00;
RAM[16'h1D7E] = 8'h00;
RAM[16'h1D7F] = 8'h00;
RAM[16'h1D80] = 8'h00;
RAM[16'h1D81] = 8'h00;
RAM[16'h1D82] = 8'h00;
RAM[16'h1D83] = 8'h00;
RAM[16'h1D84] = 8'h00;
RAM[16'h1D85] = 8'h00;
RAM[16'h1D86] = 8'h00;
RAM[16'h1D87] = 8'h00;
RAM[16'h1D88] = 8'h00;
RAM[16'h1D89] = 8'h00;
RAM[16'h1D8A] = 8'h00;
RAM[16'h1D8B] = 8'h00;
RAM[16'h1D8C] = 8'h00;
RAM[16'h1D8D] = 8'h00;
RAM[16'h1D8E] = 8'h00;
RAM[16'h1D8F] = 8'h00;
RAM[16'h1D90] = 8'h00;
RAM[16'h1D91] = 8'h00;
RAM[16'h1D92] = 8'h00;
RAM[16'h1D93] = 8'h00;
RAM[16'h1D94] = 8'h00;
RAM[16'h1D95] = 8'h00;
RAM[16'h1D96] = 8'h00;
RAM[16'h1D97] = 8'h00;
RAM[16'h1D98] = 8'h00;
RAM[16'h1D99] = 8'h00;
RAM[16'h1D9A] = 8'h00;
RAM[16'h1D9B] = 8'h00;
RAM[16'h1D9C] = 8'h00;
RAM[16'h1D9D] = 8'h00;
RAM[16'h1D9E] = 8'h00;
RAM[16'h1D9F] = 8'h00;
RAM[16'h1DA0] = 8'h00;
RAM[16'h1DA1] = 8'h00;
RAM[16'h1DA2] = 8'h00;
RAM[16'h1DA3] = 8'h00;
RAM[16'h1DA4] = 8'h00;
RAM[16'h1DA5] = 8'h00;
RAM[16'h1DA6] = 8'h00;
RAM[16'h1DA7] = 8'h00;
RAM[16'h1DA8] = 8'h00;
RAM[16'h1DA9] = 8'h00;
RAM[16'h1DAA] = 8'h00;
RAM[16'h1DAB] = 8'h00;
RAM[16'h1DAC] = 8'h00;
RAM[16'h1DAD] = 8'h00;
RAM[16'h1DAE] = 8'h00;
RAM[16'h1DAF] = 8'h00;
RAM[16'h1DB0] = 8'h00;
RAM[16'h1DB1] = 8'h00;
RAM[16'h1DB2] = 8'h00;
RAM[16'h1DB3] = 8'h00;
RAM[16'h1DB4] = 8'h00;
RAM[16'h1DB5] = 8'h00;
RAM[16'h1DB6] = 8'h00;
RAM[16'h1DB7] = 8'h00;
RAM[16'h1DB8] = 8'h00;
RAM[16'h1DB9] = 8'h00;
RAM[16'h1DBA] = 8'h00;
RAM[16'h1DBB] = 8'h00;
RAM[16'h1DBC] = 8'h00;
RAM[16'h1DBD] = 8'h00;
RAM[16'h1DBE] = 8'h00;
RAM[16'h1DBF] = 8'h00;
RAM[16'h1DC0] = 8'h00;
RAM[16'h1DC1] = 8'h00;
RAM[16'h1DC2] = 8'h00;
RAM[16'h1DC3] = 8'h00;
RAM[16'h1DC4] = 8'h00;
RAM[16'h1DC5] = 8'h00;
RAM[16'h1DC6] = 8'h00;
RAM[16'h1DC7] = 8'h00;
RAM[16'h1DC8] = 8'h00;
RAM[16'h1DC9] = 8'h00;
RAM[16'h1DCA] = 8'h00;
RAM[16'h1DCB] = 8'h00;
RAM[16'h1DCC] = 8'h00;
RAM[16'h1DCD] = 8'h00;
RAM[16'h1DCE] = 8'h00;
RAM[16'h1DCF] = 8'h00;
RAM[16'h1DD0] = 8'h00;
RAM[16'h1DD1] = 8'h00;
RAM[16'h1DD2] = 8'h00;
RAM[16'h1DD3] = 8'h00;
RAM[16'h1DD4] = 8'h00;
RAM[16'h1DD5] = 8'h00;
RAM[16'h1DD6] = 8'h00;
RAM[16'h1DD7] = 8'h00;
RAM[16'h1DD8] = 8'h00;
RAM[16'h1DD9] = 8'h00;
RAM[16'h1DDA] = 8'h00;
RAM[16'h1DDB] = 8'h00;
RAM[16'h1DDC] = 8'h00;
RAM[16'h1DDD] = 8'h00;
RAM[16'h1DDE] = 8'h00;
RAM[16'h1DDF] = 8'h00;
RAM[16'h1DE0] = 8'h00;
RAM[16'h1DE1] = 8'h00;
RAM[16'h1DE2] = 8'h00;
RAM[16'h1DE3] = 8'h00;
RAM[16'h1DE4] = 8'h00;
RAM[16'h1DE5] = 8'h00;
RAM[16'h1DE6] = 8'h00;
RAM[16'h1DE7] = 8'h00;
RAM[16'h1DE8] = 8'h00;
RAM[16'h1DE9] = 8'h00;
RAM[16'h1DEA] = 8'h00;
RAM[16'h1DEB] = 8'h00;
RAM[16'h1DEC] = 8'h00;
RAM[16'h1DED] = 8'h00;
RAM[16'h1DEE] = 8'h00;
RAM[16'h1DEF] = 8'h00;
RAM[16'h1DF0] = 8'h00;
RAM[16'h1DF1] = 8'h00;
RAM[16'h1DF2] = 8'h00;
RAM[16'h1DF3] = 8'h00;
RAM[16'h1DF4] = 8'h00;
RAM[16'h1DF5] = 8'h00;
RAM[16'h1DF6] = 8'h00;
RAM[16'h1DF7] = 8'h00;
RAM[16'h1DF8] = 8'h00;
RAM[16'h1DF9] = 8'h00;
RAM[16'h1DFA] = 8'h00;
RAM[16'h1DFB] = 8'h00;
RAM[16'h1DFC] = 8'h00;
RAM[16'h1DFD] = 8'h00;
RAM[16'h1DFE] = 8'h00;
RAM[16'h1DFF] = 8'h00;
RAM[16'h1E00] = 8'h00;
RAM[16'h1E01] = 8'h00;
RAM[16'h1E02] = 8'h00;
RAM[16'h1E03] = 8'h00;
RAM[16'h1E04] = 8'h00;
RAM[16'h1E05] = 8'h00;
RAM[16'h1E06] = 8'h00;
RAM[16'h1E07] = 8'h00;
RAM[16'h1E08] = 8'h00;
RAM[16'h1E09] = 8'h00;
RAM[16'h1E0A] = 8'h00;
RAM[16'h1E0B] = 8'h00;
RAM[16'h1E0C] = 8'h00;
RAM[16'h1E0D] = 8'h00;
RAM[16'h1E0E] = 8'h00;
RAM[16'h1E0F] = 8'h00;
RAM[16'h1E10] = 8'h00;
RAM[16'h1E11] = 8'h00;
RAM[16'h1E12] = 8'h00;
RAM[16'h1E13] = 8'h00;
RAM[16'h1E14] = 8'h00;
RAM[16'h1E15] = 8'h00;
RAM[16'h1E16] = 8'h00;
RAM[16'h1E17] = 8'h00;
RAM[16'h1E18] = 8'h00;
RAM[16'h1E19] = 8'h00;
RAM[16'h1E1A] = 8'h00;
RAM[16'h1E1B] = 8'h00;
RAM[16'h1E1C] = 8'h00;
RAM[16'h1E1D] = 8'h00;
RAM[16'h1E1E] = 8'h00;
RAM[16'h1E1F] = 8'h00;
RAM[16'h1E20] = 8'h00;
RAM[16'h1E21] = 8'h00;
RAM[16'h1E22] = 8'h00;
RAM[16'h1E23] = 8'h00;
RAM[16'h1E24] = 8'h00;
RAM[16'h1E25] = 8'h00;
RAM[16'h1E26] = 8'h00;
RAM[16'h1E27] = 8'h00;
RAM[16'h1E28] = 8'h00;
RAM[16'h1E29] = 8'h00;
RAM[16'h1E2A] = 8'h00;
RAM[16'h1E2B] = 8'h00;
RAM[16'h1E2C] = 8'h00;
RAM[16'h1E2D] = 8'h00;
RAM[16'h1E2E] = 8'h00;
RAM[16'h1E2F] = 8'h00;
RAM[16'h1E30] = 8'h00;
RAM[16'h1E31] = 8'h00;
RAM[16'h1E32] = 8'h00;
RAM[16'h1E33] = 8'h00;
RAM[16'h1E34] = 8'h00;
RAM[16'h1E35] = 8'h00;
RAM[16'h1E36] = 8'h00;
RAM[16'h1E37] = 8'h00;
RAM[16'h1E38] = 8'h00;
RAM[16'h1E39] = 8'h00;
RAM[16'h1E3A] = 8'h00;
RAM[16'h1E3B] = 8'h00;
RAM[16'h1E3C] = 8'h00;
RAM[16'h1E3D] = 8'h00;
RAM[16'h1E3E] = 8'h00;
RAM[16'h1E3F] = 8'h00;
RAM[16'h1E40] = 8'h00;
RAM[16'h1E41] = 8'h00;
RAM[16'h1E42] = 8'h00;
RAM[16'h1E43] = 8'h00;
RAM[16'h1E44] = 8'h00;
RAM[16'h1E45] = 8'h00;
RAM[16'h1E46] = 8'h00;
RAM[16'h1E47] = 8'h00;
RAM[16'h1E48] = 8'h00;
RAM[16'h1E49] = 8'h00;
RAM[16'h1E4A] = 8'h00;
RAM[16'h1E4B] = 8'h00;
RAM[16'h1E4C] = 8'h00;
RAM[16'h1E4D] = 8'h00;
RAM[16'h1E4E] = 8'h00;
RAM[16'h1E4F] = 8'h00;
RAM[16'h1E50] = 8'h00;
RAM[16'h1E51] = 8'h00;
RAM[16'h1E52] = 8'h00;
RAM[16'h1E53] = 8'h00;
RAM[16'h1E54] = 8'h00;
RAM[16'h1E55] = 8'h00;
RAM[16'h1E56] = 8'h00;
RAM[16'h1E57] = 8'h00;
RAM[16'h1E58] = 8'h00;
RAM[16'h1E59] = 8'h00;
RAM[16'h1E5A] = 8'h00;
RAM[16'h1E5B] = 8'h00;
RAM[16'h1E5C] = 8'h00;
RAM[16'h1E5D] = 8'h00;
RAM[16'h1E5E] = 8'h00;
RAM[16'h1E5F] = 8'h00;
RAM[16'h1E60] = 8'h00;
RAM[16'h1E61] = 8'h00;
RAM[16'h1E62] = 8'h00;
RAM[16'h1E63] = 8'h00;
RAM[16'h1E64] = 8'h00;
RAM[16'h1E65] = 8'h00;
RAM[16'h1E66] = 8'h00;
RAM[16'h1E67] = 8'h00;
RAM[16'h1E68] = 8'h00;
RAM[16'h1E69] = 8'h00;
RAM[16'h1E6A] = 8'h00;
RAM[16'h1E6B] = 8'h00;
RAM[16'h1E6C] = 8'h00;
RAM[16'h1E6D] = 8'h00;
RAM[16'h1E6E] = 8'h00;
RAM[16'h1E6F] = 8'h00;
RAM[16'h1E70] = 8'h00;
RAM[16'h1E71] = 8'h00;
RAM[16'h1E72] = 8'h00;
RAM[16'h1E73] = 8'h00;
RAM[16'h1E74] = 8'h00;
RAM[16'h1E75] = 8'h00;
RAM[16'h1E76] = 8'h00;
RAM[16'h1E77] = 8'h00;
RAM[16'h1E78] = 8'h00;
RAM[16'h1E79] = 8'h00;
RAM[16'h1E7A] = 8'h00;
RAM[16'h1E7B] = 8'h00;
RAM[16'h1E7C] = 8'h00;
RAM[16'h1E7D] = 8'h00;
RAM[16'h1E7E] = 8'h00;
RAM[16'h1E7F] = 8'h00;
RAM[16'h1E80] = 8'h00;
RAM[16'h1E81] = 8'h00;
RAM[16'h1E82] = 8'h00;
RAM[16'h1E83] = 8'h00;
RAM[16'h1E84] = 8'h00;
RAM[16'h1E85] = 8'h00;
RAM[16'h1E86] = 8'h00;
RAM[16'h1E87] = 8'h00;
RAM[16'h1E88] = 8'h00;
RAM[16'h1E89] = 8'h00;
RAM[16'h1E8A] = 8'h00;
RAM[16'h1E8B] = 8'h00;
RAM[16'h1E8C] = 8'h00;
RAM[16'h1E8D] = 8'h00;
RAM[16'h1E8E] = 8'h00;
RAM[16'h1E8F] = 8'h00;
RAM[16'h1E90] = 8'h00;
RAM[16'h1E91] = 8'h00;
RAM[16'h1E92] = 8'h00;
RAM[16'h1E93] = 8'h00;
RAM[16'h1E94] = 8'h00;
RAM[16'h1E95] = 8'h00;
RAM[16'h1E96] = 8'h00;
RAM[16'h1E97] = 8'h00;
RAM[16'h1E98] = 8'h00;
RAM[16'h1E99] = 8'h00;
RAM[16'h1E9A] = 8'h00;
RAM[16'h1E9B] = 8'h00;
RAM[16'h1E9C] = 8'h00;
RAM[16'h1E9D] = 8'h00;
RAM[16'h1E9E] = 8'h00;
RAM[16'h1E9F] = 8'h00;
RAM[16'h1EA0] = 8'h00;
RAM[16'h1EA1] = 8'h00;
RAM[16'h1EA2] = 8'h00;
RAM[16'h1EA3] = 8'h00;
RAM[16'h1EA4] = 8'h00;
RAM[16'h1EA5] = 8'h00;
RAM[16'h1EA6] = 8'h00;
RAM[16'h1EA7] = 8'h00;
RAM[16'h1EA8] = 8'h00;
RAM[16'h1EA9] = 8'h00;
RAM[16'h1EAA] = 8'h00;
RAM[16'h1EAB] = 8'h00;
RAM[16'h1EAC] = 8'h00;
RAM[16'h1EAD] = 8'h00;
RAM[16'h1EAE] = 8'h00;
RAM[16'h1EAF] = 8'h00;
RAM[16'h1EB0] = 8'h00;
RAM[16'h1EB1] = 8'h00;
RAM[16'h1EB2] = 8'h00;
RAM[16'h1EB3] = 8'h00;
RAM[16'h1EB4] = 8'h00;
RAM[16'h1EB5] = 8'h00;
RAM[16'h1EB6] = 8'h00;
RAM[16'h1EB7] = 8'h00;
RAM[16'h1EB8] = 8'h00;
RAM[16'h1EB9] = 8'h00;
RAM[16'h1EBA] = 8'h00;
RAM[16'h1EBB] = 8'h00;
RAM[16'h1EBC] = 8'h00;
RAM[16'h1EBD] = 8'h00;
RAM[16'h1EBE] = 8'h00;
RAM[16'h1EBF] = 8'h00;
RAM[16'h1EC0] = 8'h00;
RAM[16'h1EC1] = 8'h00;
RAM[16'h1EC2] = 8'h00;
RAM[16'h1EC3] = 8'h00;
RAM[16'h1EC4] = 8'h00;
RAM[16'h1EC5] = 8'h00;
RAM[16'h1EC6] = 8'h00;
RAM[16'h1EC7] = 8'h00;
RAM[16'h1EC8] = 8'h00;
RAM[16'h1EC9] = 8'h00;
RAM[16'h1ECA] = 8'h00;
RAM[16'h1ECB] = 8'h00;
RAM[16'h1ECC] = 8'h00;
RAM[16'h1ECD] = 8'h00;
RAM[16'h1ECE] = 8'h00;
RAM[16'h1ECF] = 8'h00;
RAM[16'h1ED0] = 8'h00;
RAM[16'h1ED1] = 8'h00;
RAM[16'h1ED2] = 8'h00;
RAM[16'h1ED3] = 8'h00;
RAM[16'h1ED4] = 8'h00;
RAM[16'h1ED5] = 8'h00;
RAM[16'h1ED6] = 8'h00;
RAM[16'h1ED7] = 8'h00;
RAM[16'h1ED8] = 8'h00;
RAM[16'h1ED9] = 8'h00;
RAM[16'h1EDA] = 8'h00;
RAM[16'h1EDB] = 8'h00;
RAM[16'h1EDC] = 8'h00;
RAM[16'h1EDD] = 8'h00;
RAM[16'h1EDE] = 8'h00;
RAM[16'h1EDF] = 8'h00;
RAM[16'h1EE0] = 8'h00;
RAM[16'h1EE1] = 8'h00;
RAM[16'h1EE2] = 8'h00;
RAM[16'h1EE3] = 8'h00;
RAM[16'h1EE4] = 8'h00;
RAM[16'h1EE5] = 8'h00;
RAM[16'h1EE6] = 8'h00;
RAM[16'h1EE7] = 8'h00;
RAM[16'h1EE8] = 8'h00;
RAM[16'h1EE9] = 8'h00;
RAM[16'h1EEA] = 8'h00;
RAM[16'h1EEB] = 8'h00;
RAM[16'h1EEC] = 8'h00;
RAM[16'h1EED] = 8'h00;
RAM[16'h1EEE] = 8'h00;
RAM[16'h1EEF] = 8'h00;
RAM[16'h1EF0] = 8'h00;
RAM[16'h1EF1] = 8'h00;
RAM[16'h1EF2] = 8'h00;
RAM[16'h1EF3] = 8'h00;
RAM[16'h1EF4] = 8'h00;
RAM[16'h1EF5] = 8'h00;
RAM[16'h1EF6] = 8'h00;
RAM[16'h1EF7] = 8'h00;
RAM[16'h1EF8] = 8'h00;
RAM[16'h1EF9] = 8'h00;
RAM[16'h1EFA] = 8'h00;
RAM[16'h1EFB] = 8'h00;
RAM[16'h1EFC] = 8'h00;
RAM[16'h1EFD] = 8'h00;
RAM[16'h1EFE] = 8'h00;
RAM[16'h1EFF] = 8'h00;
RAM[16'h1F00] = 8'h00;
RAM[16'h1F01] = 8'h00;
RAM[16'h1F02] = 8'h00;
RAM[16'h1F03] = 8'h00;
RAM[16'h1F04] = 8'h00;
RAM[16'h1F05] = 8'h00;
RAM[16'h1F06] = 8'h00;
RAM[16'h1F07] = 8'h00;
RAM[16'h1F08] = 8'h00;
RAM[16'h1F09] = 8'h00;
RAM[16'h1F0A] = 8'h00;
RAM[16'h1F0B] = 8'h00;
RAM[16'h1F0C] = 8'h00;
RAM[16'h1F0D] = 8'h00;
RAM[16'h1F0E] = 8'h00;
RAM[16'h1F0F] = 8'h00;
RAM[16'h1F10] = 8'h00;
RAM[16'h1F11] = 8'h00;
RAM[16'h1F12] = 8'h00;
RAM[16'h1F13] = 8'h00;
RAM[16'h1F14] = 8'h00;
RAM[16'h1F15] = 8'h00;
RAM[16'h1F16] = 8'h00;
RAM[16'h1F17] = 8'h00;
RAM[16'h1F18] = 8'h00;
RAM[16'h1F19] = 8'h00;
RAM[16'h1F1A] = 8'h00;
RAM[16'h1F1B] = 8'h00;
RAM[16'h1F1C] = 8'h00;
RAM[16'h1F1D] = 8'h00;
RAM[16'h1F1E] = 8'h00;
RAM[16'h1F1F] = 8'h00;
RAM[16'h1F20] = 8'h00;
RAM[16'h1F21] = 8'h00;
RAM[16'h1F22] = 8'h00;
RAM[16'h1F23] = 8'h00;
RAM[16'h1F24] = 8'h00;
RAM[16'h1F25] = 8'h00;
RAM[16'h1F26] = 8'h00;
RAM[16'h1F27] = 8'h00;
RAM[16'h1F28] = 8'h00;
RAM[16'h1F29] = 8'h00;
RAM[16'h1F2A] = 8'h00;
RAM[16'h1F2B] = 8'h00;
RAM[16'h1F2C] = 8'h00;
RAM[16'h1F2D] = 8'h00;
RAM[16'h1F2E] = 8'h00;
RAM[16'h1F2F] = 8'h00;
RAM[16'h1F30] = 8'h00;
RAM[16'h1F31] = 8'h00;
RAM[16'h1F32] = 8'h00;
RAM[16'h1F33] = 8'h00;
RAM[16'h1F34] = 8'h00;
RAM[16'h1F35] = 8'h00;
RAM[16'h1F36] = 8'h00;
RAM[16'h1F37] = 8'h00;
RAM[16'h1F38] = 8'h00;
RAM[16'h1F39] = 8'h00;
RAM[16'h1F3A] = 8'h00;
RAM[16'h1F3B] = 8'h00;
RAM[16'h1F3C] = 8'h00;
RAM[16'h1F3D] = 8'h00;
RAM[16'h1F3E] = 8'h00;
RAM[16'h1F3F] = 8'h00;
RAM[16'h1F40] = 8'h00;
RAM[16'h1F41] = 8'h00;
RAM[16'h1F42] = 8'h00;
RAM[16'h1F43] = 8'h00;
RAM[16'h1F44] = 8'h00;
RAM[16'h1F45] = 8'h00;
RAM[16'h1F46] = 8'h00;
RAM[16'h1F47] = 8'h00;
RAM[16'h1F48] = 8'h00;
RAM[16'h1F49] = 8'h00;
RAM[16'h1F4A] = 8'h00;
RAM[16'h1F4B] = 8'h00;
RAM[16'h1F4C] = 8'h00;
RAM[16'h1F4D] = 8'h00;
RAM[16'h1F4E] = 8'h00;
RAM[16'h1F4F] = 8'h00;
RAM[16'h1F50] = 8'h00;
RAM[16'h1F51] = 8'h00;
RAM[16'h1F52] = 8'h00;
RAM[16'h1F53] = 8'h00;
RAM[16'h1F54] = 8'h00;
RAM[16'h1F55] = 8'h00;
RAM[16'h1F56] = 8'h00;
RAM[16'h1F57] = 8'h00;
RAM[16'h1F58] = 8'h00;
RAM[16'h1F59] = 8'h00;
RAM[16'h1F5A] = 8'h00;
RAM[16'h1F5B] = 8'h00;
RAM[16'h1F5C] = 8'h00;
RAM[16'h1F5D] = 8'h00;
RAM[16'h1F5E] = 8'h00;
RAM[16'h1F5F] = 8'h00;
RAM[16'h1F60] = 8'h00;
RAM[16'h1F61] = 8'h00;
RAM[16'h1F62] = 8'h00;
RAM[16'h1F63] = 8'h00;
RAM[16'h1F64] = 8'h00;
RAM[16'h1F65] = 8'h00;
RAM[16'h1F66] = 8'h00;
RAM[16'h1F67] = 8'h00;
RAM[16'h1F68] = 8'h00;
RAM[16'h1F69] = 8'h00;
RAM[16'h1F6A] = 8'h00;
RAM[16'h1F6B] = 8'h00;
RAM[16'h1F6C] = 8'h00;
RAM[16'h1F6D] = 8'h00;
RAM[16'h1F6E] = 8'h00;
RAM[16'h1F6F] = 8'h00;
RAM[16'h1F70] = 8'h00;
RAM[16'h1F71] = 8'h00;
RAM[16'h1F72] = 8'h00;
RAM[16'h1F73] = 8'h00;
RAM[16'h1F74] = 8'h00;
RAM[16'h1F75] = 8'h00;
RAM[16'h1F76] = 8'h00;
RAM[16'h1F77] = 8'h00;
RAM[16'h1F78] = 8'h00;
RAM[16'h1F79] = 8'h00;
RAM[16'h1F7A] = 8'h00;
RAM[16'h1F7B] = 8'h00;
RAM[16'h1F7C] = 8'h00;
RAM[16'h1F7D] = 8'h00;
RAM[16'h1F7E] = 8'h00;
RAM[16'h1F7F] = 8'h00;
RAM[16'h1F80] = 8'h00;
RAM[16'h1F81] = 8'h00;
RAM[16'h1F82] = 8'h00;
RAM[16'h1F83] = 8'h00;
RAM[16'h1F84] = 8'h00;
RAM[16'h1F85] = 8'h00;
RAM[16'h1F86] = 8'h00;
RAM[16'h1F87] = 8'h00;
RAM[16'h1F88] = 8'h00;
RAM[16'h1F89] = 8'h00;
RAM[16'h1F8A] = 8'h00;
RAM[16'h1F8B] = 8'h00;
RAM[16'h1F8C] = 8'h00;
RAM[16'h1F8D] = 8'h00;
RAM[16'h1F8E] = 8'h00;
RAM[16'h1F8F] = 8'h00;
RAM[16'h1F90] = 8'h00;
RAM[16'h1F91] = 8'h00;
RAM[16'h1F92] = 8'h00;
RAM[16'h1F93] = 8'h00;
RAM[16'h1F94] = 8'h00;
RAM[16'h1F95] = 8'h00;
RAM[16'h1F96] = 8'h00;
RAM[16'h1F97] = 8'h00;
RAM[16'h1F98] = 8'h00;
RAM[16'h1F99] = 8'h00;
RAM[16'h1F9A] = 8'h00;
RAM[16'h1F9B] = 8'h00;
RAM[16'h1F9C] = 8'h00;
RAM[16'h1F9D] = 8'h00;
RAM[16'h1F9E] = 8'h00;
RAM[16'h1F9F] = 8'h00;
RAM[16'h1FA0] = 8'h00;
RAM[16'h1FA1] = 8'h00;
RAM[16'h1FA2] = 8'h00;
RAM[16'h1FA3] = 8'h00;
RAM[16'h1FA4] = 8'h00;
RAM[16'h1FA5] = 8'h00;
RAM[16'h1FA6] = 8'h00;
RAM[16'h1FA7] = 8'h00;
RAM[16'h1FA8] = 8'h00;
RAM[16'h1FA9] = 8'h00;
RAM[16'h1FAA] = 8'h00;
RAM[16'h1FAB] = 8'h00;
RAM[16'h1FAC] = 8'h00;
RAM[16'h1FAD] = 8'h00;
RAM[16'h1FAE] = 8'h00;
RAM[16'h1FAF] = 8'h00;
RAM[16'h1FB0] = 8'h00;
RAM[16'h1FB1] = 8'h00;
RAM[16'h1FB2] = 8'h00;
RAM[16'h1FB3] = 8'h00;
RAM[16'h1FB4] = 8'h00;
RAM[16'h1FB5] = 8'h00;
RAM[16'h1FB6] = 8'h00;
RAM[16'h1FB7] = 8'h00;
RAM[16'h1FB8] = 8'h00;
RAM[16'h1FB9] = 8'h00;
RAM[16'h1FBA] = 8'h00;
RAM[16'h1FBB] = 8'h00;
RAM[16'h1FBC] = 8'h00;
RAM[16'h1FBD] = 8'h00;
RAM[16'h1FBE] = 8'h00;
RAM[16'h1FBF] = 8'h00;
RAM[16'h1FC0] = 8'h00;
RAM[16'h1FC1] = 8'h00;
RAM[16'h1FC2] = 8'h00;
RAM[16'h1FC3] = 8'h00;
RAM[16'h1FC4] = 8'h00;
RAM[16'h1FC5] = 8'h00;
RAM[16'h1FC6] = 8'h00;
RAM[16'h1FC7] = 8'h00;
RAM[16'h1FC8] = 8'h00;
RAM[16'h1FC9] = 8'h00;
RAM[16'h1FCA] = 8'h00;
RAM[16'h1FCB] = 8'h00;
RAM[16'h1FCC] = 8'h00;
RAM[16'h1FCD] = 8'h00;
RAM[16'h1FCE] = 8'h00;
RAM[16'h1FCF] = 8'h00;
RAM[16'h1FD0] = 8'h00;
RAM[16'h1FD1] = 8'h00;
RAM[16'h1FD2] = 8'h00;
RAM[16'h1FD3] = 8'h00;
RAM[16'h1FD4] = 8'h00;
RAM[16'h1FD5] = 8'h00;
RAM[16'h1FD6] = 8'h00;
RAM[16'h1FD7] = 8'h00;
RAM[16'h1FD8] = 8'h00;
RAM[16'h1FD9] = 8'h00;
RAM[16'h1FDA] = 8'h00;
RAM[16'h1FDB] = 8'h00;
RAM[16'h1FDC] = 8'h00;
RAM[16'h1FDD] = 8'h00;
RAM[16'h1FDE] = 8'h00;
RAM[16'h1FDF] = 8'h00;
RAM[16'h1FE0] = 8'h00;
RAM[16'h1FE1] = 8'h00;
RAM[16'h1FE2] = 8'h00;
RAM[16'h1FE3] = 8'h00;
RAM[16'h1FE4] = 8'h00;
RAM[16'h1FE5] = 8'h00;
RAM[16'h1FE6] = 8'h00;
RAM[16'h1FE7] = 8'h00;
RAM[16'h1FE8] = 8'h00;
RAM[16'h1FE9] = 8'h00;
RAM[16'h1FEA] = 8'h00;
RAM[16'h1FEB] = 8'h00;
RAM[16'h1FEC] = 8'h00;
RAM[16'h1FED] = 8'h00;
RAM[16'h1FEE] = 8'h00;
RAM[16'h1FEF] = 8'h00;
RAM[16'h1FF0] = 8'h00;
RAM[16'h1FF1] = 8'h00;
RAM[16'h1FF2] = 8'h00;
RAM[16'h1FF3] = 8'h00;
RAM[16'h1FF4] = 8'h00;
RAM[16'h1FF5] = 8'h00;
RAM[16'h1FF6] = 8'h00;
RAM[16'h1FF7] = 8'h00;
RAM[16'h1FF8] = 8'h00;
RAM[16'h1FF9] = 8'h00;
RAM[16'h1FFA] = 8'h00;
RAM[16'h1FFB] = 8'h00;
RAM[16'h1FFC] = 8'h00;
RAM[16'h1FFD] = 8'h00;
RAM[16'h1FFE] = 8'h00;
RAM[16'h1FFF] = 8'h00;
RAM[16'h2000] = 8'h00;
RAM[16'h2001] = 8'h00;
RAM[16'h2002] = 8'h00;
RAM[16'h2003] = 8'h00;
RAM[16'h2004] = 8'h00;
RAM[16'h2005] = 8'h00;
RAM[16'h2006] = 8'h00;
RAM[16'h2007] = 8'h00;
RAM[16'h2008] = 8'h00;
RAM[16'h2009] = 8'h00;
RAM[16'h200A] = 8'h00;
RAM[16'h200B] = 8'h00;
RAM[16'h200C] = 8'h00;
RAM[16'h200D] = 8'h00;
RAM[16'h200E] = 8'h00;
RAM[16'h200F] = 8'h00;
RAM[16'h2010] = 8'h00;
RAM[16'h2011] = 8'h00;
RAM[16'h2012] = 8'h00;
RAM[16'h2013] = 8'h00;
RAM[16'h2014] = 8'h00;
RAM[16'h2015] = 8'h00;
RAM[16'h2016] = 8'h00;
RAM[16'h2017] = 8'h00;
RAM[16'h2018] = 8'h00;
RAM[16'h2019] = 8'h00;
RAM[16'h201A] = 8'h00;
RAM[16'h201B] = 8'h00;
RAM[16'h201C] = 8'h00;
RAM[16'h201D] = 8'h00;
RAM[16'h201E] = 8'h00;
RAM[16'h201F] = 8'h00;
RAM[16'h2020] = 8'h00;
RAM[16'h2021] = 8'h00;
RAM[16'h2022] = 8'h00;
RAM[16'h2023] = 8'h00;
RAM[16'h2024] = 8'h00;
RAM[16'h2025] = 8'h00;
RAM[16'h2026] = 8'h00;
RAM[16'h2027] = 8'h00;
RAM[16'h2028] = 8'h00;
RAM[16'h2029] = 8'h00;
RAM[16'h202A] = 8'h00;
RAM[16'h202B] = 8'h00;
RAM[16'h202C] = 8'h00;
RAM[16'h202D] = 8'h00;
RAM[16'h202E] = 8'h00;
RAM[16'h202F] = 8'h00;
RAM[16'h2030] = 8'h00;
RAM[16'h2031] = 8'h00;
RAM[16'h2032] = 8'h00;
RAM[16'h2033] = 8'h00;
RAM[16'h2034] = 8'h00;
RAM[16'h2035] = 8'h00;
RAM[16'h2036] = 8'h00;
RAM[16'h2037] = 8'h00;
RAM[16'h2038] = 8'h00;
RAM[16'h2039] = 8'h00;
RAM[16'h203A] = 8'h00;
RAM[16'h203B] = 8'h00;
RAM[16'h203C] = 8'h00;
RAM[16'h203D] = 8'h00;
RAM[16'h203E] = 8'h00;
RAM[16'h203F] = 8'h00;
RAM[16'h2040] = 8'h00;
RAM[16'h2041] = 8'h00;
RAM[16'h2042] = 8'h00;
RAM[16'h2043] = 8'h00;
RAM[16'h2044] = 8'h00;
RAM[16'h2045] = 8'h00;
RAM[16'h2046] = 8'h00;
RAM[16'h2047] = 8'h00;
RAM[16'h2048] = 8'h00;
RAM[16'h2049] = 8'h00;
RAM[16'h204A] = 8'h00;
RAM[16'h204B] = 8'h00;
RAM[16'h204C] = 8'h00;
RAM[16'h204D] = 8'h00;
RAM[16'h204E] = 8'h00;
RAM[16'h204F] = 8'h00;
RAM[16'h2050] = 8'h00;
RAM[16'h2051] = 8'h00;
RAM[16'h2052] = 8'h00;
RAM[16'h2053] = 8'h00;
RAM[16'h2054] = 8'h00;
RAM[16'h2055] = 8'h00;
RAM[16'h2056] = 8'h00;
RAM[16'h2057] = 8'h00;
RAM[16'h2058] = 8'h00;
RAM[16'h2059] = 8'h00;
RAM[16'h205A] = 8'h00;
RAM[16'h205B] = 8'h00;
RAM[16'h205C] = 8'h00;
RAM[16'h205D] = 8'h00;
RAM[16'h205E] = 8'h00;
RAM[16'h205F] = 8'h00;
RAM[16'h2060] = 8'h00;
RAM[16'h2061] = 8'h00;
RAM[16'h2062] = 8'h00;
RAM[16'h2063] = 8'h00;
RAM[16'h2064] = 8'h00;
RAM[16'h2065] = 8'h00;
RAM[16'h2066] = 8'h00;
RAM[16'h2067] = 8'h00;
RAM[16'h2068] = 8'h00;
RAM[16'h2069] = 8'h00;
RAM[16'h206A] = 8'h00;
RAM[16'h206B] = 8'h00;
RAM[16'h206C] = 8'h00;
RAM[16'h206D] = 8'h00;
RAM[16'h206E] = 8'h00;
RAM[16'h206F] = 8'h00;
RAM[16'h2070] = 8'h00;
RAM[16'h2071] = 8'h00;
RAM[16'h2072] = 8'h00;
RAM[16'h2073] = 8'h00;
RAM[16'h2074] = 8'h00;
RAM[16'h2075] = 8'h00;
RAM[16'h2076] = 8'h00;
RAM[16'h2077] = 8'h00;
RAM[16'h2078] = 8'h00;
RAM[16'h2079] = 8'h00;
RAM[16'h207A] = 8'h00;
RAM[16'h207B] = 8'h00;
RAM[16'h207C] = 8'h00;
RAM[16'h207D] = 8'h00;
RAM[16'h207E] = 8'h00;
RAM[16'h207F] = 8'h00;
RAM[16'h2080] = 8'h00;
RAM[16'h2081] = 8'h00;
RAM[16'h2082] = 8'h00;
RAM[16'h2083] = 8'h00;
RAM[16'h2084] = 8'h00;
RAM[16'h2085] = 8'h00;
RAM[16'h2086] = 8'h00;
RAM[16'h2087] = 8'h00;
RAM[16'h2088] = 8'h00;
RAM[16'h2089] = 8'h00;
RAM[16'h208A] = 8'h00;
RAM[16'h208B] = 8'h00;
RAM[16'h208C] = 8'h00;
RAM[16'h208D] = 8'h00;
RAM[16'h208E] = 8'h00;
RAM[16'h208F] = 8'h00;
RAM[16'h2090] = 8'h00;
RAM[16'h2091] = 8'h00;
RAM[16'h2092] = 8'h00;
RAM[16'h2093] = 8'h00;
RAM[16'h2094] = 8'h00;
RAM[16'h2095] = 8'h00;
RAM[16'h2096] = 8'h00;
RAM[16'h2097] = 8'h00;
RAM[16'h2098] = 8'h00;
RAM[16'h2099] = 8'h00;
RAM[16'h209A] = 8'h00;
RAM[16'h209B] = 8'h00;
RAM[16'h209C] = 8'h00;
RAM[16'h209D] = 8'h00;
RAM[16'h209E] = 8'h00;
RAM[16'h209F] = 8'h00;
RAM[16'h20A0] = 8'h00;
RAM[16'h20A1] = 8'h00;
RAM[16'h20A2] = 8'h00;
RAM[16'h20A3] = 8'h00;
RAM[16'h20A4] = 8'h00;
RAM[16'h20A5] = 8'h00;
RAM[16'h20A6] = 8'h00;
RAM[16'h20A7] = 8'h00;
RAM[16'h20A8] = 8'h00;
RAM[16'h20A9] = 8'h00;
RAM[16'h20AA] = 8'h00;
RAM[16'h20AB] = 8'h00;
RAM[16'h20AC] = 8'h00;
RAM[16'h20AD] = 8'h00;
RAM[16'h20AE] = 8'h00;
RAM[16'h20AF] = 8'h00;
RAM[16'h20B0] = 8'h00;
RAM[16'h20B1] = 8'h00;
RAM[16'h20B2] = 8'h00;
RAM[16'h20B3] = 8'h00;
RAM[16'h20B4] = 8'h00;
RAM[16'h20B5] = 8'h00;
RAM[16'h20B6] = 8'h00;
RAM[16'h20B7] = 8'h00;
RAM[16'h20B8] = 8'h00;
RAM[16'h20B9] = 8'h00;
RAM[16'h20BA] = 8'h00;
RAM[16'h20BB] = 8'h00;
RAM[16'h20BC] = 8'h00;
RAM[16'h20BD] = 8'h00;
RAM[16'h20BE] = 8'h00;
RAM[16'h20BF] = 8'h00;
RAM[16'h20C0] = 8'h00;
RAM[16'h20C1] = 8'h00;
RAM[16'h20C2] = 8'h00;
RAM[16'h20C3] = 8'h00;
RAM[16'h20C4] = 8'h00;
RAM[16'h20C5] = 8'h00;
RAM[16'h20C6] = 8'h00;
RAM[16'h20C7] = 8'h00;
RAM[16'h20C8] = 8'h00;
RAM[16'h20C9] = 8'h00;
RAM[16'h20CA] = 8'h00;
RAM[16'h20CB] = 8'h00;
RAM[16'h20CC] = 8'h00;
RAM[16'h20CD] = 8'h00;
RAM[16'h20CE] = 8'h00;
RAM[16'h20CF] = 8'h00;
RAM[16'h20D0] = 8'h00;
RAM[16'h20D1] = 8'h00;
RAM[16'h20D2] = 8'h00;
RAM[16'h20D3] = 8'h00;
RAM[16'h20D4] = 8'h00;
RAM[16'h20D5] = 8'h00;
RAM[16'h20D6] = 8'h00;
RAM[16'h20D7] = 8'h00;
RAM[16'h20D8] = 8'h00;
RAM[16'h20D9] = 8'h00;
RAM[16'h20DA] = 8'h00;
RAM[16'h20DB] = 8'h00;
RAM[16'h20DC] = 8'h00;
RAM[16'h20DD] = 8'h00;
RAM[16'h20DE] = 8'h00;
RAM[16'h20DF] = 8'h00;
RAM[16'h20E0] = 8'h00;
RAM[16'h20E1] = 8'h00;
RAM[16'h20E2] = 8'h00;
RAM[16'h20E3] = 8'h00;
RAM[16'h20E4] = 8'h00;
RAM[16'h20E5] = 8'h00;
RAM[16'h20E6] = 8'h00;
RAM[16'h20E7] = 8'h00;
RAM[16'h20E8] = 8'h00;
RAM[16'h20E9] = 8'h00;
RAM[16'h20EA] = 8'h00;
RAM[16'h20EB] = 8'h00;
RAM[16'h20EC] = 8'h00;
RAM[16'h20ED] = 8'h00;
RAM[16'h20EE] = 8'h00;
RAM[16'h20EF] = 8'h00;
RAM[16'h20F0] = 8'h00;
RAM[16'h20F1] = 8'h00;
RAM[16'h20F2] = 8'h00;
RAM[16'h20F3] = 8'h00;
RAM[16'h20F4] = 8'h00;
RAM[16'h20F5] = 8'h00;
RAM[16'h20F6] = 8'h00;
RAM[16'h20F7] = 8'h00;
RAM[16'h20F8] = 8'h00;
RAM[16'h20F9] = 8'h00;
RAM[16'h20FA] = 8'h00;
RAM[16'h20FB] = 8'h00;
RAM[16'h20FC] = 8'h00;
RAM[16'h20FD] = 8'h00;
RAM[16'h20FE] = 8'h00;
RAM[16'h20FF] = 8'h00;
RAM[16'h2100] = 8'h00;
RAM[16'h2101] = 8'h00;
RAM[16'h2102] = 8'h00;
RAM[16'h2103] = 8'h00;
RAM[16'h2104] = 8'h00;
RAM[16'h2105] = 8'h00;
RAM[16'h2106] = 8'h00;
RAM[16'h2107] = 8'h00;
RAM[16'h2108] = 8'h00;
RAM[16'h2109] = 8'h00;
RAM[16'h210A] = 8'h00;
RAM[16'h210B] = 8'h00;
RAM[16'h210C] = 8'h00;
RAM[16'h210D] = 8'h00;
RAM[16'h210E] = 8'h00;
RAM[16'h210F] = 8'h00;
RAM[16'h2110] = 8'h00;
RAM[16'h2111] = 8'h00;
RAM[16'h2112] = 8'h00;
RAM[16'h2113] = 8'h00;
RAM[16'h2114] = 8'h00;
RAM[16'h2115] = 8'h00;
RAM[16'h2116] = 8'h00;
RAM[16'h2117] = 8'h00;
RAM[16'h2118] = 8'h00;
RAM[16'h2119] = 8'h00;
RAM[16'h211A] = 8'h00;
RAM[16'h211B] = 8'h00;
RAM[16'h211C] = 8'h00;
RAM[16'h211D] = 8'h00;
RAM[16'h211E] = 8'h00;
RAM[16'h211F] = 8'h00;
RAM[16'h2120] = 8'h00;
RAM[16'h2121] = 8'h00;
RAM[16'h2122] = 8'h00;
RAM[16'h2123] = 8'h00;
RAM[16'h2124] = 8'h00;
RAM[16'h2125] = 8'h00;
RAM[16'h2126] = 8'h00;
RAM[16'h2127] = 8'h00;
RAM[16'h2128] = 8'h00;
RAM[16'h2129] = 8'h00;
RAM[16'h212A] = 8'h00;
RAM[16'h212B] = 8'h00;
RAM[16'h212C] = 8'h00;
RAM[16'h212D] = 8'h00;
RAM[16'h212E] = 8'h00;
RAM[16'h212F] = 8'h00;
RAM[16'h2130] = 8'h00;
RAM[16'h2131] = 8'h00;
RAM[16'h2132] = 8'h00;
RAM[16'h2133] = 8'h00;
RAM[16'h2134] = 8'h00;
RAM[16'h2135] = 8'h00;
RAM[16'h2136] = 8'h00;
RAM[16'h2137] = 8'h00;
RAM[16'h2138] = 8'h00;
RAM[16'h2139] = 8'h00;
RAM[16'h213A] = 8'h00;
RAM[16'h213B] = 8'h00;
RAM[16'h213C] = 8'h00;
RAM[16'h213D] = 8'h00;
RAM[16'h213E] = 8'h00;
RAM[16'h213F] = 8'h00;
RAM[16'h2140] = 8'h00;
RAM[16'h2141] = 8'h00;
RAM[16'h2142] = 8'h00;
RAM[16'h2143] = 8'h00;
RAM[16'h2144] = 8'h00;
RAM[16'h2145] = 8'h00;
RAM[16'h2146] = 8'h00;
RAM[16'h2147] = 8'h00;
RAM[16'h2148] = 8'h00;
RAM[16'h2149] = 8'h00;
RAM[16'h214A] = 8'h00;
RAM[16'h214B] = 8'h00;
RAM[16'h214C] = 8'h00;
RAM[16'h214D] = 8'h00;
RAM[16'h214E] = 8'h00;
RAM[16'h214F] = 8'h00;
RAM[16'h2150] = 8'h00;
RAM[16'h2151] = 8'h00;
RAM[16'h2152] = 8'h00;
RAM[16'h2153] = 8'h00;
RAM[16'h2154] = 8'h00;
RAM[16'h2155] = 8'h00;
RAM[16'h2156] = 8'h00;
RAM[16'h2157] = 8'h00;
RAM[16'h2158] = 8'h00;
RAM[16'h2159] = 8'h00;
RAM[16'h215A] = 8'h00;
RAM[16'h215B] = 8'h00;
RAM[16'h215C] = 8'h00;
RAM[16'h215D] = 8'h00;
RAM[16'h215E] = 8'h00;
RAM[16'h215F] = 8'h00;
RAM[16'h2160] = 8'h00;
RAM[16'h2161] = 8'h00;
RAM[16'h2162] = 8'h00;
RAM[16'h2163] = 8'h00;
RAM[16'h2164] = 8'h00;
RAM[16'h2165] = 8'h00;
RAM[16'h2166] = 8'h00;
RAM[16'h2167] = 8'h00;
RAM[16'h2168] = 8'h00;
RAM[16'h2169] = 8'h00;
RAM[16'h216A] = 8'h00;
RAM[16'h216B] = 8'h00;
RAM[16'h216C] = 8'h00;
RAM[16'h216D] = 8'h00;
RAM[16'h216E] = 8'h00;
RAM[16'h216F] = 8'h00;
RAM[16'h2170] = 8'h00;
RAM[16'h2171] = 8'h00;
RAM[16'h2172] = 8'h00;
RAM[16'h2173] = 8'h00;
RAM[16'h2174] = 8'h00;
RAM[16'h2175] = 8'h00;
RAM[16'h2176] = 8'h00;
RAM[16'h2177] = 8'h00;
RAM[16'h2178] = 8'h00;
RAM[16'h2179] = 8'h00;
RAM[16'h217A] = 8'h00;
RAM[16'h217B] = 8'h00;
RAM[16'h217C] = 8'h00;
RAM[16'h217D] = 8'h00;
RAM[16'h217E] = 8'h00;
RAM[16'h217F] = 8'h00;
RAM[16'h2180] = 8'h00;
RAM[16'h2181] = 8'h00;
RAM[16'h2182] = 8'h00;
RAM[16'h2183] = 8'h00;
RAM[16'h2184] = 8'h00;
RAM[16'h2185] = 8'h00;
RAM[16'h2186] = 8'h00;
RAM[16'h2187] = 8'h00;
RAM[16'h2188] = 8'h00;
RAM[16'h2189] = 8'h00;
RAM[16'h218A] = 8'h00;
RAM[16'h218B] = 8'h00;
RAM[16'h218C] = 8'h00;
RAM[16'h218D] = 8'h00;
RAM[16'h218E] = 8'h00;
RAM[16'h218F] = 8'h00;
RAM[16'h2190] = 8'h00;
RAM[16'h2191] = 8'h00;
RAM[16'h2192] = 8'h00;
RAM[16'h2193] = 8'h00;
RAM[16'h2194] = 8'h00;
RAM[16'h2195] = 8'h00;
RAM[16'h2196] = 8'h00;
RAM[16'h2197] = 8'h00;
RAM[16'h2198] = 8'h00;
RAM[16'h2199] = 8'h00;
RAM[16'h219A] = 8'h00;
RAM[16'h219B] = 8'h00;
RAM[16'h219C] = 8'h00;
RAM[16'h219D] = 8'h00;
RAM[16'h219E] = 8'h00;
RAM[16'h219F] = 8'h00;
RAM[16'h21A0] = 8'h00;
RAM[16'h21A1] = 8'h00;
RAM[16'h21A2] = 8'h00;
RAM[16'h21A3] = 8'h00;
RAM[16'h21A4] = 8'h00;
RAM[16'h21A5] = 8'h00;
RAM[16'h21A6] = 8'h00;
RAM[16'h21A7] = 8'h00;
RAM[16'h21A8] = 8'h00;
RAM[16'h21A9] = 8'h00;
RAM[16'h21AA] = 8'h00;
RAM[16'h21AB] = 8'h00;
RAM[16'h21AC] = 8'h00;
RAM[16'h21AD] = 8'h00;
RAM[16'h21AE] = 8'h00;
RAM[16'h21AF] = 8'h00;
RAM[16'h21B0] = 8'h00;
RAM[16'h21B1] = 8'h00;
RAM[16'h21B2] = 8'h00;
RAM[16'h21B3] = 8'h00;
RAM[16'h21B4] = 8'h00;
RAM[16'h21B5] = 8'h00;
RAM[16'h21B6] = 8'h00;
RAM[16'h21B7] = 8'h00;
RAM[16'h21B8] = 8'h00;
RAM[16'h21B9] = 8'h00;
RAM[16'h21BA] = 8'h00;
RAM[16'h21BB] = 8'h00;
RAM[16'h21BC] = 8'h00;
RAM[16'h21BD] = 8'h00;
RAM[16'h21BE] = 8'h00;
RAM[16'h21BF] = 8'h00;
RAM[16'h21C0] = 8'h00;
RAM[16'h21C1] = 8'h00;
RAM[16'h21C2] = 8'h00;
RAM[16'h21C3] = 8'h00;
RAM[16'h21C4] = 8'h00;
RAM[16'h21C5] = 8'h00;
RAM[16'h21C6] = 8'h00;
RAM[16'h21C7] = 8'h00;
RAM[16'h21C8] = 8'h00;
RAM[16'h21C9] = 8'h00;
RAM[16'h21CA] = 8'h00;
RAM[16'h21CB] = 8'h00;
RAM[16'h21CC] = 8'h00;
RAM[16'h21CD] = 8'h00;
RAM[16'h21CE] = 8'h00;
RAM[16'h21CF] = 8'h00;
RAM[16'h21D0] = 8'h00;
RAM[16'h21D1] = 8'h00;
RAM[16'h21D2] = 8'h00;
RAM[16'h21D3] = 8'h00;
RAM[16'h21D4] = 8'h00;
RAM[16'h21D5] = 8'h00;
RAM[16'h21D6] = 8'h00;
RAM[16'h21D7] = 8'h00;
RAM[16'h21D8] = 8'h00;
RAM[16'h21D9] = 8'h00;
RAM[16'h21DA] = 8'h00;
RAM[16'h21DB] = 8'h00;
RAM[16'h21DC] = 8'h00;
RAM[16'h21DD] = 8'h00;
RAM[16'h21DE] = 8'h00;
RAM[16'h21DF] = 8'h00;
RAM[16'h21E0] = 8'h00;
RAM[16'h21E1] = 8'h00;
RAM[16'h21E2] = 8'h00;
RAM[16'h21E3] = 8'h00;
RAM[16'h21E4] = 8'h00;
RAM[16'h21E5] = 8'h00;
RAM[16'h21E6] = 8'h00;
RAM[16'h21E7] = 8'h00;
RAM[16'h21E8] = 8'h00;
RAM[16'h21E9] = 8'h00;
RAM[16'h21EA] = 8'h00;
RAM[16'h21EB] = 8'h00;
RAM[16'h21EC] = 8'h00;
RAM[16'h21ED] = 8'h00;
RAM[16'h21EE] = 8'h00;
RAM[16'h21EF] = 8'h00;
RAM[16'h21F0] = 8'h00;
RAM[16'h21F1] = 8'h00;
RAM[16'h21F2] = 8'h00;
RAM[16'h21F3] = 8'h00;
RAM[16'h21F4] = 8'h00;
RAM[16'h21F5] = 8'h00;
RAM[16'h21F6] = 8'h00;
RAM[16'h21F7] = 8'h00;
RAM[16'h21F8] = 8'h00;
RAM[16'h21F9] = 8'h00;
RAM[16'h21FA] = 8'h00;
RAM[16'h21FB] = 8'h00;
RAM[16'h21FC] = 8'h00;
RAM[16'h21FD] = 8'h00;
RAM[16'h21FE] = 8'h00;
RAM[16'h21FF] = 8'h00;
RAM[16'h2200] = 8'h00;
RAM[16'h2201] = 8'h00;
RAM[16'h2202] = 8'h00;
RAM[16'h2203] = 8'h00;
RAM[16'h2204] = 8'h00;
RAM[16'h2205] = 8'h00;
RAM[16'h2206] = 8'h00;
RAM[16'h2207] = 8'h00;
RAM[16'h2208] = 8'h00;
RAM[16'h2209] = 8'h00;
RAM[16'h220A] = 8'h00;
RAM[16'h220B] = 8'h00;
RAM[16'h220C] = 8'h00;
RAM[16'h220D] = 8'h00;
RAM[16'h220E] = 8'h00;
RAM[16'h220F] = 8'h00;
RAM[16'h2210] = 8'h00;
RAM[16'h2211] = 8'h00;
RAM[16'h2212] = 8'h00;
RAM[16'h2213] = 8'h00;
RAM[16'h2214] = 8'h00;
RAM[16'h2215] = 8'h00;
RAM[16'h2216] = 8'h00;
RAM[16'h2217] = 8'h00;
RAM[16'h2218] = 8'h00;
RAM[16'h2219] = 8'h00;
RAM[16'h221A] = 8'h00;
RAM[16'h221B] = 8'h00;
RAM[16'h221C] = 8'h00;
RAM[16'h221D] = 8'h00;
RAM[16'h221E] = 8'h00;
RAM[16'h221F] = 8'h00;
RAM[16'h2220] = 8'h00;
RAM[16'h2221] = 8'h00;
RAM[16'h2222] = 8'h00;
RAM[16'h2223] = 8'h00;
RAM[16'h2224] = 8'h00;
RAM[16'h2225] = 8'h00;
RAM[16'h2226] = 8'h00;
RAM[16'h2227] = 8'h00;
RAM[16'h2228] = 8'h00;
RAM[16'h2229] = 8'h00;
RAM[16'h222A] = 8'h00;
RAM[16'h222B] = 8'h00;
RAM[16'h222C] = 8'h00;
RAM[16'h222D] = 8'h00;
RAM[16'h222E] = 8'h00;
RAM[16'h222F] = 8'h00;
RAM[16'h2230] = 8'h00;
RAM[16'h2231] = 8'h00;
RAM[16'h2232] = 8'h00;
RAM[16'h2233] = 8'h00;
RAM[16'h2234] = 8'h00;
RAM[16'h2235] = 8'h00;
RAM[16'h2236] = 8'h00;
RAM[16'h2237] = 8'h00;
RAM[16'h2238] = 8'h00;
RAM[16'h2239] = 8'h00;
RAM[16'h223A] = 8'h00;
RAM[16'h223B] = 8'h00;
RAM[16'h223C] = 8'h00;
RAM[16'h223D] = 8'h00;
RAM[16'h223E] = 8'h00;
RAM[16'h223F] = 8'h00;
RAM[16'h2240] = 8'h00;
RAM[16'h2241] = 8'h00;
RAM[16'h2242] = 8'h00;
RAM[16'h2243] = 8'h00;
RAM[16'h2244] = 8'h00;
RAM[16'h2245] = 8'h00;
RAM[16'h2246] = 8'h00;
RAM[16'h2247] = 8'h00;
RAM[16'h2248] = 8'h00;
RAM[16'h2249] = 8'h00;
RAM[16'h224A] = 8'h00;
RAM[16'h224B] = 8'h00;
RAM[16'h224C] = 8'h00;
RAM[16'h224D] = 8'h00;
RAM[16'h224E] = 8'h00;
RAM[16'h224F] = 8'h00;
RAM[16'h2250] = 8'h00;
RAM[16'h2251] = 8'h00;
RAM[16'h2252] = 8'h00;
RAM[16'h2253] = 8'h00;
RAM[16'h2254] = 8'h00;
RAM[16'h2255] = 8'h00;
RAM[16'h2256] = 8'h00;
RAM[16'h2257] = 8'h00;
RAM[16'h2258] = 8'h00;
RAM[16'h2259] = 8'h00;
RAM[16'h225A] = 8'h00;
RAM[16'h225B] = 8'h00;
RAM[16'h225C] = 8'h00;
RAM[16'h225D] = 8'h00;
RAM[16'h225E] = 8'h00;
RAM[16'h225F] = 8'h00;
RAM[16'h2260] = 8'h00;
RAM[16'h2261] = 8'h00;
RAM[16'h2262] = 8'h00;
RAM[16'h2263] = 8'h00;
RAM[16'h2264] = 8'h00;
RAM[16'h2265] = 8'h00;
RAM[16'h2266] = 8'h00;
RAM[16'h2267] = 8'h00;
RAM[16'h2268] = 8'h00;
RAM[16'h2269] = 8'h00;
RAM[16'h226A] = 8'h00;
RAM[16'h226B] = 8'h00;
RAM[16'h226C] = 8'h00;
RAM[16'h226D] = 8'h00;
RAM[16'h226E] = 8'h00;
RAM[16'h226F] = 8'h00;
RAM[16'h2270] = 8'h00;
RAM[16'h2271] = 8'h00;
RAM[16'h2272] = 8'h00;
RAM[16'h2273] = 8'h00;
RAM[16'h2274] = 8'h00;
RAM[16'h2275] = 8'h00;
RAM[16'h2276] = 8'h00;
RAM[16'h2277] = 8'h00;
RAM[16'h2278] = 8'h00;
RAM[16'h2279] = 8'h00;
RAM[16'h227A] = 8'h00;
RAM[16'h227B] = 8'h00;
RAM[16'h227C] = 8'h00;
RAM[16'h227D] = 8'h00;
RAM[16'h227E] = 8'h00;
RAM[16'h227F] = 8'h00;
RAM[16'h2280] = 8'h00;
RAM[16'h2281] = 8'h00;
RAM[16'h2282] = 8'h00;
RAM[16'h2283] = 8'h00;
RAM[16'h2284] = 8'h00;
RAM[16'h2285] = 8'h00;
RAM[16'h2286] = 8'h00;
RAM[16'h2287] = 8'h00;
RAM[16'h2288] = 8'h00;
RAM[16'h2289] = 8'h00;
RAM[16'h228A] = 8'h00;
RAM[16'h228B] = 8'h00;
RAM[16'h228C] = 8'h00;
RAM[16'h228D] = 8'h00;
RAM[16'h228E] = 8'h00;
RAM[16'h228F] = 8'h00;
RAM[16'h2290] = 8'h00;
RAM[16'h2291] = 8'h00;
RAM[16'h2292] = 8'h00;
RAM[16'h2293] = 8'h00;
RAM[16'h2294] = 8'h00;
RAM[16'h2295] = 8'h00;
RAM[16'h2296] = 8'h00;
RAM[16'h2297] = 8'h00;
RAM[16'h2298] = 8'h00;
RAM[16'h2299] = 8'h00;
RAM[16'h229A] = 8'h00;
RAM[16'h229B] = 8'h00;
RAM[16'h229C] = 8'h00;
RAM[16'h229D] = 8'h00;
RAM[16'h229E] = 8'h00;
RAM[16'h229F] = 8'h00;
RAM[16'h22A0] = 8'h00;
RAM[16'h22A1] = 8'h00;
RAM[16'h22A2] = 8'h00;
RAM[16'h22A3] = 8'h00;
RAM[16'h22A4] = 8'h00;
RAM[16'h22A5] = 8'h00;
RAM[16'h22A6] = 8'h00;
RAM[16'h22A7] = 8'h00;
RAM[16'h22A8] = 8'h00;
RAM[16'h22A9] = 8'h00;
RAM[16'h22AA] = 8'h00;
RAM[16'h22AB] = 8'h00;
RAM[16'h22AC] = 8'h00;
RAM[16'h22AD] = 8'h00;
RAM[16'h22AE] = 8'h00;
RAM[16'h22AF] = 8'h00;
RAM[16'h22B0] = 8'h00;
RAM[16'h22B1] = 8'h00;
RAM[16'h22B2] = 8'h00;
RAM[16'h22B3] = 8'h00;
RAM[16'h22B4] = 8'h00;
RAM[16'h22B5] = 8'h00;
RAM[16'h22B6] = 8'h00;
RAM[16'h22B7] = 8'h00;
RAM[16'h22B8] = 8'h00;
RAM[16'h22B9] = 8'h00;
RAM[16'h22BA] = 8'h00;
RAM[16'h22BB] = 8'h00;
RAM[16'h22BC] = 8'h00;
RAM[16'h22BD] = 8'h00;
RAM[16'h22BE] = 8'h00;
RAM[16'h22BF] = 8'h00;
RAM[16'h22C0] = 8'h00;
RAM[16'h22C1] = 8'h00;
RAM[16'h22C2] = 8'h00;
RAM[16'h22C3] = 8'h00;
RAM[16'h22C4] = 8'h00;
RAM[16'h22C5] = 8'h00;
RAM[16'h22C6] = 8'h00;
RAM[16'h22C7] = 8'h00;
RAM[16'h22C8] = 8'h00;
RAM[16'h22C9] = 8'h00;
RAM[16'h22CA] = 8'h00;
RAM[16'h22CB] = 8'h00;
RAM[16'h22CC] = 8'h00;
RAM[16'h22CD] = 8'h00;
RAM[16'h22CE] = 8'h00;
RAM[16'h22CF] = 8'h00;
RAM[16'h22D0] = 8'h00;
RAM[16'h22D1] = 8'h00;
RAM[16'h22D2] = 8'h00;
RAM[16'h22D3] = 8'h00;
RAM[16'h22D4] = 8'h00;
RAM[16'h22D5] = 8'h00;
RAM[16'h22D6] = 8'h00;
RAM[16'h22D7] = 8'h00;
RAM[16'h22D8] = 8'h00;
RAM[16'h22D9] = 8'h00;
RAM[16'h22DA] = 8'h00;
RAM[16'h22DB] = 8'h00;
RAM[16'h22DC] = 8'h00;
RAM[16'h22DD] = 8'h00;
RAM[16'h22DE] = 8'h00;
RAM[16'h22DF] = 8'h00;
RAM[16'h22E0] = 8'h00;
RAM[16'h22E1] = 8'h00;
RAM[16'h22E2] = 8'h00;
RAM[16'h22E3] = 8'h00;
RAM[16'h22E4] = 8'h00;
RAM[16'h22E5] = 8'h00;
RAM[16'h22E6] = 8'h00;
RAM[16'h22E7] = 8'h00;
RAM[16'h22E8] = 8'h00;
RAM[16'h22E9] = 8'h00;
RAM[16'h22EA] = 8'h00;
RAM[16'h22EB] = 8'h00;
RAM[16'h22EC] = 8'h00;
RAM[16'h22ED] = 8'h00;
RAM[16'h22EE] = 8'h00;
RAM[16'h22EF] = 8'h00;
RAM[16'h22F0] = 8'h00;
RAM[16'h22F1] = 8'h00;
RAM[16'h22F2] = 8'h00;
RAM[16'h22F3] = 8'h00;
RAM[16'h22F4] = 8'h00;
RAM[16'h22F5] = 8'h00;
RAM[16'h22F6] = 8'h00;
RAM[16'h22F7] = 8'h00;
RAM[16'h22F8] = 8'h00;
RAM[16'h22F9] = 8'h00;
RAM[16'h22FA] = 8'h00;
RAM[16'h22FB] = 8'h00;
RAM[16'h22FC] = 8'h00;
RAM[16'h22FD] = 8'h00;
RAM[16'h22FE] = 8'h00;
RAM[16'h22FF] = 8'h00;
RAM[16'h2300] = 8'h00;
RAM[16'h2301] = 8'h00;
RAM[16'h2302] = 8'h00;
RAM[16'h2303] = 8'h00;
RAM[16'h2304] = 8'h00;
RAM[16'h2305] = 8'h00;
RAM[16'h2306] = 8'h00;
RAM[16'h2307] = 8'h00;
RAM[16'h2308] = 8'h00;
RAM[16'h2309] = 8'h00;
RAM[16'h230A] = 8'h00;
RAM[16'h230B] = 8'h00;
RAM[16'h230C] = 8'h00;
RAM[16'h230D] = 8'h00;
RAM[16'h230E] = 8'h00;
RAM[16'h230F] = 8'h00;
RAM[16'h2310] = 8'h00;
RAM[16'h2311] = 8'h00;
RAM[16'h2312] = 8'h00;
RAM[16'h2313] = 8'h00;
RAM[16'h2314] = 8'h00;
RAM[16'h2315] = 8'h00;
RAM[16'h2316] = 8'h00;
RAM[16'h2317] = 8'h00;
RAM[16'h2318] = 8'h00;
RAM[16'h2319] = 8'h00;
RAM[16'h231A] = 8'h00;
RAM[16'h231B] = 8'h00;
RAM[16'h231C] = 8'h00;
RAM[16'h231D] = 8'h00;
RAM[16'h231E] = 8'h00;
RAM[16'h231F] = 8'h00;
RAM[16'h2320] = 8'h00;
RAM[16'h2321] = 8'h00;
RAM[16'h2322] = 8'h00;
RAM[16'h2323] = 8'h00;
RAM[16'h2324] = 8'h00;
RAM[16'h2325] = 8'h00;
RAM[16'h2326] = 8'h00;
RAM[16'h2327] = 8'h00;
RAM[16'h2328] = 8'h00;
RAM[16'h2329] = 8'h00;
RAM[16'h232A] = 8'h00;
RAM[16'h232B] = 8'h00;
RAM[16'h232C] = 8'h00;
RAM[16'h232D] = 8'h00;
RAM[16'h232E] = 8'h00;
RAM[16'h232F] = 8'h00;
RAM[16'h2330] = 8'h00;
RAM[16'h2331] = 8'h00;
RAM[16'h2332] = 8'h00;
RAM[16'h2333] = 8'h00;
RAM[16'h2334] = 8'h00;
RAM[16'h2335] = 8'h00;
RAM[16'h2336] = 8'h00;
RAM[16'h2337] = 8'h00;
RAM[16'h2338] = 8'h00;
RAM[16'h2339] = 8'h00;
RAM[16'h233A] = 8'h00;
RAM[16'h233B] = 8'h00;
RAM[16'h233C] = 8'h00;
RAM[16'h233D] = 8'h00;
RAM[16'h233E] = 8'h00;
RAM[16'h233F] = 8'h00;
RAM[16'h2340] = 8'h00;
RAM[16'h2341] = 8'h00;
RAM[16'h2342] = 8'h00;
RAM[16'h2343] = 8'h00;
RAM[16'h2344] = 8'h00;
RAM[16'h2345] = 8'h00;
RAM[16'h2346] = 8'h00;
RAM[16'h2347] = 8'h00;
RAM[16'h2348] = 8'h00;
RAM[16'h2349] = 8'h00;
RAM[16'h234A] = 8'h00;
RAM[16'h234B] = 8'h00;
RAM[16'h234C] = 8'h00;
RAM[16'h234D] = 8'h00;
RAM[16'h234E] = 8'h00;
RAM[16'h234F] = 8'h00;
RAM[16'h2350] = 8'h00;
RAM[16'h2351] = 8'h00;
RAM[16'h2352] = 8'h00;
RAM[16'h2353] = 8'h00;
RAM[16'h2354] = 8'h00;
RAM[16'h2355] = 8'h00;
RAM[16'h2356] = 8'h00;
RAM[16'h2357] = 8'h00;
RAM[16'h2358] = 8'h00;
RAM[16'h2359] = 8'h00;
RAM[16'h235A] = 8'h00;
RAM[16'h235B] = 8'h00;
RAM[16'h235C] = 8'h00;
RAM[16'h235D] = 8'h00;
RAM[16'h235E] = 8'h00;
RAM[16'h235F] = 8'h00;
RAM[16'h2360] = 8'h00;
RAM[16'h2361] = 8'h00;
RAM[16'h2362] = 8'h00;
RAM[16'h2363] = 8'h00;
RAM[16'h2364] = 8'h00;
RAM[16'h2365] = 8'h00;
RAM[16'h2366] = 8'h00;
RAM[16'h2367] = 8'h00;
RAM[16'h2368] = 8'h00;
RAM[16'h2369] = 8'h00;
RAM[16'h236A] = 8'h00;
RAM[16'h236B] = 8'h00;
RAM[16'h236C] = 8'h00;
RAM[16'h236D] = 8'h00;
RAM[16'h236E] = 8'h00;
RAM[16'h236F] = 8'h00;
RAM[16'h2370] = 8'h00;
RAM[16'h2371] = 8'h00;
RAM[16'h2372] = 8'h00;
RAM[16'h2373] = 8'h00;
RAM[16'h2374] = 8'h00;
RAM[16'h2375] = 8'h00;
RAM[16'h2376] = 8'h00;
RAM[16'h2377] = 8'h00;
RAM[16'h2378] = 8'h00;
RAM[16'h2379] = 8'h00;
RAM[16'h237A] = 8'h00;
RAM[16'h237B] = 8'h00;
RAM[16'h237C] = 8'h00;
RAM[16'h237D] = 8'h00;
RAM[16'h237E] = 8'h00;
RAM[16'h237F] = 8'h00;
RAM[16'h2380] = 8'h00;
RAM[16'h2381] = 8'h00;
RAM[16'h2382] = 8'h00;
RAM[16'h2383] = 8'h00;
RAM[16'h2384] = 8'h00;
RAM[16'h2385] = 8'h00;
RAM[16'h2386] = 8'h00;
RAM[16'h2387] = 8'h00;
RAM[16'h2388] = 8'h00;
RAM[16'h2389] = 8'h00;
RAM[16'h238A] = 8'h00;
RAM[16'h238B] = 8'h00;
RAM[16'h238C] = 8'h00;
RAM[16'h238D] = 8'h00;
RAM[16'h238E] = 8'h00;
RAM[16'h238F] = 8'h00;
RAM[16'h2390] = 8'h00;
RAM[16'h2391] = 8'h00;
RAM[16'h2392] = 8'h00;
RAM[16'h2393] = 8'h00;
RAM[16'h2394] = 8'h00;
RAM[16'h2395] = 8'h00;
RAM[16'h2396] = 8'h00;
RAM[16'h2397] = 8'h00;
RAM[16'h2398] = 8'h00;
RAM[16'h2399] = 8'h00;
RAM[16'h239A] = 8'h00;
RAM[16'h239B] = 8'h00;
RAM[16'h239C] = 8'h00;
RAM[16'h239D] = 8'h00;
RAM[16'h239E] = 8'h00;
RAM[16'h239F] = 8'h00;
RAM[16'h23A0] = 8'h00;
RAM[16'h23A1] = 8'h00;
RAM[16'h23A2] = 8'h00;
RAM[16'h23A3] = 8'h00;
RAM[16'h23A4] = 8'h00;
RAM[16'h23A5] = 8'h00;
RAM[16'h23A6] = 8'h00;
RAM[16'h23A7] = 8'h00;
RAM[16'h23A8] = 8'h00;
RAM[16'h23A9] = 8'h00;
RAM[16'h23AA] = 8'h00;
RAM[16'h23AB] = 8'h00;
RAM[16'h23AC] = 8'h00;
RAM[16'h23AD] = 8'h00;
RAM[16'h23AE] = 8'h00;
RAM[16'h23AF] = 8'h00;
RAM[16'h23B0] = 8'h00;
RAM[16'h23B1] = 8'h00;
RAM[16'h23B2] = 8'h00;
RAM[16'h23B3] = 8'h00;
RAM[16'h23B4] = 8'h00;
RAM[16'h23B5] = 8'h00;
RAM[16'h23B6] = 8'h00;
RAM[16'h23B7] = 8'h00;
RAM[16'h23B8] = 8'h00;
RAM[16'h23B9] = 8'h00;
RAM[16'h23BA] = 8'h00;
RAM[16'h23BB] = 8'h00;
RAM[16'h23BC] = 8'h00;
RAM[16'h23BD] = 8'h00;
RAM[16'h23BE] = 8'h00;
RAM[16'h23BF] = 8'h00;
RAM[16'h23C0] = 8'h00;
RAM[16'h23C1] = 8'h00;
RAM[16'h23C2] = 8'h00;
RAM[16'h23C3] = 8'h00;
RAM[16'h23C4] = 8'h00;
RAM[16'h23C5] = 8'h00;
RAM[16'h23C6] = 8'h00;
RAM[16'h23C7] = 8'h00;
RAM[16'h23C8] = 8'h00;
RAM[16'h23C9] = 8'h00;
RAM[16'h23CA] = 8'h00;
RAM[16'h23CB] = 8'h00;
RAM[16'h23CC] = 8'h00;
RAM[16'h23CD] = 8'h00;
RAM[16'h23CE] = 8'h00;
RAM[16'h23CF] = 8'h00;
RAM[16'h23D0] = 8'h00;
RAM[16'h23D1] = 8'h00;
RAM[16'h23D2] = 8'h00;
RAM[16'h23D3] = 8'h00;
RAM[16'h23D4] = 8'h00;
RAM[16'h23D5] = 8'h00;
RAM[16'h23D6] = 8'h00;
RAM[16'h23D7] = 8'h00;
RAM[16'h23D8] = 8'h00;
RAM[16'h23D9] = 8'h00;
RAM[16'h23DA] = 8'h00;
RAM[16'h23DB] = 8'h00;
RAM[16'h23DC] = 8'h00;
RAM[16'h23DD] = 8'h00;
RAM[16'h23DE] = 8'h00;
RAM[16'h23DF] = 8'h00;
RAM[16'h23E0] = 8'h00;
RAM[16'h23E1] = 8'h00;
RAM[16'h23E2] = 8'h00;
RAM[16'h23E3] = 8'h00;
RAM[16'h23E4] = 8'h00;
RAM[16'h23E5] = 8'h00;
RAM[16'h23E6] = 8'h00;
RAM[16'h23E7] = 8'h00;
RAM[16'h23E8] = 8'h00;
RAM[16'h23E9] = 8'h00;
RAM[16'h23EA] = 8'h00;
RAM[16'h23EB] = 8'h00;
RAM[16'h23EC] = 8'h00;
RAM[16'h23ED] = 8'h00;
RAM[16'h23EE] = 8'h00;
RAM[16'h23EF] = 8'h00;
RAM[16'h23F0] = 8'h00;
RAM[16'h23F1] = 8'h00;
RAM[16'h23F2] = 8'h00;
RAM[16'h23F3] = 8'h00;
RAM[16'h23F4] = 8'h00;
RAM[16'h23F5] = 8'h00;
RAM[16'h23F6] = 8'h00;
RAM[16'h23F7] = 8'h00;
RAM[16'h23F8] = 8'h00;
RAM[16'h23F9] = 8'h00;
RAM[16'h23FA] = 8'h00;
RAM[16'h23FB] = 8'h00;
RAM[16'h23FC] = 8'h00;
RAM[16'h23FD] = 8'h00;
RAM[16'h23FE] = 8'h00;
RAM[16'h23FF] = 8'h00;
RAM[16'h2400] = 8'h00;
RAM[16'h2401] = 8'h00;
RAM[16'h2402] = 8'h00;
RAM[16'h2403] = 8'h00;
RAM[16'h2404] = 8'h00;
RAM[16'h2405] = 8'h00;
RAM[16'h2406] = 8'h00;
RAM[16'h2407] = 8'h00;
RAM[16'h2408] = 8'h00;
RAM[16'h2409] = 8'h00;
RAM[16'h240A] = 8'h00;
RAM[16'h240B] = 8'h00;
RAM[16'h240C] = 8'h00;
RAM[16'h240D] = 8'h00;
RAM[16'h240E] = 8'h00;
RAM[16'h240F] = 8'h00;
RAM[16'h2410] = 8'h00;
RAM[16'h2411] = 8'h00;
RAM[16'h2412] = 8'h00;
RAM[16'h2413] = 8'h00;
RAM[16'h2414] = 8'h00;
RAM[16'h2415] = 8'h00;
RAM[16'h2416] = 8'h00;
RAM[16'h2417] = 8'h00;
RAM[16'h2418] = 8'h00;
RAM[16'h2419] = 8'h00;
RAM[16'h241A] = 8'h00;
RAM[16'h241B] = 8'h00;
RAM[16'h241C] = 8'h00;
RAM[16'h241D] = 8'h00;
RAM[16'h241E] = 8'h00;
RAM[16'h241F] = 8'h00;
RAM[16'h2420] = 8'h00;
RAM[16'h2421] = 8'h00;
RAM[16'h2422] = 8'h00;
RAM[16'h2423] = 8'h00;
RAM[16'h2424] = 8'h00;
RAM[16'h2425] = 8'h00;
RAM[16'h2426] = 8'h00;
RAM[16'h2427] = 8'h00;
RAM[16'h2428] = 8'h00;
RAM[16'h2429] = 8'h00;
RAM[16'h242A] = 8'h00;
RAM[16'h242B] = 8'h00;
RAM[16'h242C] = 8'h00;
RAM[16'h242D] = 8'h00;
RAM[16'h242E] = 8'h00;
RAM[16'h242F] = 8'h00;
RAM[16'h2430] = 8'h00;
RAM[16'h2431] = 8'h00;
RAM[16'h2432] = 8'h00;
RAM[16'h2433] = 8'h00;
RAM[16'h2434] = 8'h00;
RAM[16'h2435] = 8'h00;
RAM[16'h2436] = 8'h00;
RAM[16'h2437] = 8'h00;
RAM[16'h2438] = 8'h00;
RAM[16'h2439] = 8'h00;
RAM[16'h243A] = 8'h00;
RAM[16'h243B] = 8'h00;
RAM[16'h243C] = 8'h00;
RAM[16'h243D] = 8'h00;
RAM[16'h243E] = 8'h00;
RAM[16'h243F] = 8'h00;
RAM[16'h2440] = 8'h00;
RAM[16'h2441] = 8'h00;
RAM[16'h2442] = 8'h00;
RAM[16'h2443] = 8'h00;
RAM[16'h2444] = 8'h00;
RAM[16'h2445] = 8'h00;
RAM[16'h2446] = 8'h00;
RAM[16'h2447] = 8'h00;
RAM[16'h2448] = 8'h00;
RAM[16'h2449] = 8'h00;
RAM[16'h244A] = 8'h00;
RAM[16'h244B] = 8'h00;
RAM[16'h244C] = 8'h00;
RAM[16'h244D] = 8'h00;
RAM[16'h244E] = 8'h00;
RAM[16'h244F] = 8'h00;
RAM[16'h2450] = 8'h00;
RAM[16'h2451] = 8'h00;
RAM[16'h2452] = 8'h00;
RAM[16'h2453] = 8'h00;
RAM[16'h2454] = 8'h00;
RAM[16'h2455] = 8'h00;
RAM[16'h2456] = 8'h00;
RAM[16'h2457] = 8'h00;
RAM[16'h2458] = 8'h00;
RAM[16'h2459] = 8'h00;
RAM[16'h245A] = 8'h00;
RAM[16'h245B] = 8'h00;
RAM[16'h245C] = 8'h00;
RAM[16'h245D] = 8'h00;
RAM[16'h245E] = 8'h00;
RAM[16'h245F] = 8'h00;
RAM[16'h2460] = 8'h00;
RAM[16'h2461] = 8'h00;
RAM[16'h2462] = 8'h00;
RAM[16'h2463] = 8'h00;
RAM[16'h2464] = 8'h00;
RAM[16'h2465] = 8'h00;
RAM[16'h2466] = 8'h00;
RAM[16'h2467] = 8'h00;
RAM[16'h2468] = 8'h00;
RAM[16'h2469] = 8'h00;
RAM[16'h246A] = 8'h00;
RAM[16'h246B] = 8'h00;
RAM[16'h246C] = 8'h00;
RAM[16'h246D] = 8'h00;
RAM[16'h246E] = 8'h00;
RAM[16'h246F] = 8'h00;
RAM[16'h2470] = 8'h00;
RAM[16'h2471] = 8'h00;
RAM[16'h2472] = 8'h00;
RAM[16'h2473] = 8'h00;
RAM[16'h2474] = 8'h00;
RAM[16'h2475] = 8'h00;
RAM[16'h2476] = 8'h00;
RAM[16'h2477] = 8'h00;
RAM[16'h2478] = 8'h00;
RAM[16'h2479] = 8'h00;
RAM[16'h247A] = 8'h00;
RAM[16'h247B] = 8'h00;
RAM[16'h247C] = 8'h00;
RAM[16'h247D] = 8'h00;
RAM[16'h247E] = 8'h00;
RAM[16'h247F] = 8'h00;
RAM[16'h2480] = 8'h00;
RAM[16'h2481] = 8'h00;
RAM[16'h2482] = 8'h00;
RAM[16'h2483] = 8'h00;
RAM[16'h2484] = 8'h00;
RAM[16'h2485] = 8'h00;
RAM[16'h2486] = 8'h00;
RAM[16'h2487] = 8'h00;
RAM[16'h2488] = 8'h00;
RAM[16'h2489] = 8'h00;
RAM[16'h248A] = 8'h00;
RAM[16'h248B] = 8'h00;
RAM[16'h248C] = 8'h00;
RAM[16'h248D] = 8'h00;
RAM[16'h248E] = 8'h00;
RAM[16'h248F] = 8'h00;
RAM[16'h2490] = 8'h00;
RAM[16'h2491] = 8'h00;
RAM[16'h2492] = 8'h00;
RAM[16'h2493] = 8'h00;
RAM[16'h2494] = 8'h00;
RAM[16'h2495] = 8'h00;
RAM[16'h2496] = 8'h00;
RAM[16'h2497] = 8'h00;
RAM[16'h2498] = 8'h00;
RAM[16'h2499] = 8'h00;
RAM[16'h249A] = 8'h00;
RAM[16'h249B] = 8'h00;
RAM[16'h249C] = 8'h00;
RAM[16'h249D] = 8'h00;
RAM[16'h249E] = 8'h00;
RAM[16'h249F] = 8'h00;
RAM[16'h24A0] = 8'h00;
RAM[16'h24A1] = 8'h00;
RAM[16'h24A2] = 8'h00;
RAM[16'h24A3] = 8'h00;
RAM[16'h24A4] = 8'h00;
RAM[16'h24A5] = 8'h00;
RAM[16'h24A6] = 8'h00;
RAM[16'h24A7] = 8'h00;
RAM[16'h24A8] = 8'h00;
RAM[16'h24A9] = 8'h00;
RAM[16'h24AA] = 8'h00;
RAM[16'h24AB] = 8'h00;
RAM[16'h24AC] = 8'h00;
RAM[16'h24AD] = 8'h00;
RAM[16'h24AE] = 8'h00;
RAM[16'h24AF] = 8'h00;
RAM[16'h24B0] = 8'h00;
RAM[16'h24B1] = 8'h00;
RAM[16'h24B2] = 8'h00;
RAM[16'h24B3] = 8'h00;
RAM[16'h24B4] = 8'h00;
RAM[16'h24B5] = 8'h00;
RAM[16'h24B6] = 8'h00;
RAM[16'h24B7] = 8'h00;
RAM[16'h24B8] = 8'h00;
RAM[16'h24B9] = 8'h00;
RAM[16'h24BA] = 8'h00;
RAM[16'h24BB] = 8'h00;
RAM[16'h24BC] = 8'h00;
RAM[16'h24BD] = 8'h00;
RAM[16'h24BE] = 8'h00;
RAM[16'h24BF] = 8'h00;
RAM[16'h24C0] = 8'h00;
RAM[16'h24C1] = 8'h00;
RAM[16'h24C2] = 8'h00;
RAM[16'h24C3] = 8'h00;
RAM[16'h24C4] = 8'h00;
RAM[16'h24C5] = 8'h00;
RAM[16'h24C6] = 8'h00;
RAM[16'h24C7] = 8'h00;
RAM[16'h24C8] = 8'h00;
RAM[16'h24C9] = 8'h00;
RAM[16'h24CA] = 8'h00;
RAM[16'h24CB] = 8'h00;
RAM[16'h24CC] = 8'h00;
RAM[16'h24CD] = 8'h00;
RAM[16'h24CE] = 8'h00;
RAM[16'h24CF] = 8'h00;
RAM[16'h24D0] = 8'h00;
RAM[16'h24D1] = 8'h00;
RAM[16'h24D2] = 8'h00;
RAM[16'h24D3] = 8'h00;
RAM[16'h24D4] = 8'h00;
RAM[16'h24D5] = 8'h00;
RAM[16'h24D6] = 8'h00;
RAM[16'h24D7] = 8'h00;
RAM[16'h24D8] = 8'h00;
RAM[16'h24D9] = 8'h00;
RAM[16'h24DA] = 8'h00;
RAM[16'h24DB] = 8'h00;
RAM[16'h24DC] = 8'h00;
RAM[16'h24DD] = 8'h00;
RAM[16'h24DE] = 8'h00;
RAM[16'h24DF] = 8'h00;
RAM[16'h24E0] = 8'h00;
RAM[16'h24E1] = 8'h00;
RAM[16'h24E2] = 8'h00;
RAM[16'h24E3] = 8'h00;
RAM[16'h24E4] = 8'h00;
RAM[16'h24E5] = 8'h00;
RAM[16'h24E6] = 8'h00;
RAM[16'h24E7] = 8'h00;
RAM[16'h24E8] = 8'h00;
RAM[16'h24E9] = 8'h00;
RAM[16'h24EA] = 8'h00;
RAM[16'h24EB] = 8'h00;
RAM[16'h24EC] = 8'h00;
RAM[16'h24ED] = 8'h00;
RAM[16'h24EE] = 8'h00;
RAM[16'h24EF] = 8'h00;
RAM[16'h24F0] = 8'h00;
RAM[16'h24F1] = 8'h00;
RAM[16'h24F2] = 8'h00;
RAM[16'h24F3] = 8'h00;
RAM[16'h24F4] = 8'h00;
RAM[16'h24F5] = 8'h00;
RAM[16'h24F6] = 8'h00;
RAM[16'h24F7] = 8'h00;
RAM[16'h24F8] = 8'h00;
RAM[16'h24F9] = 8'h00;
RAM[16'h24FA] = 8'h00;
RAM[16'h24FB] = 8'h00;
RAM[16'h24FC] = 8'h00;
RAM[16'h24FD] = 8'h00;
RAM[16'h24FE] = 8'h00;
RAM[16'h24FF] = 8'h00;
RAM[16'h2500] = 8'h00;
RAM[16'h2501] = 8'h00;
RAM[16'h2502] = 8'h00;
RAM[16'h2503] = 8'h00;
RAM[16'h2504] = 8'h00;
RAM[16'h2505] = 8'h00;
RAM[16'h2506] = 8'h00;
RAM[16'h2507] = 8'h00;
RAM[16'h2508] = 8'h00;
RAM[16'h2509] = 8'h00;
RAM[16'h250A] = 8'h00;
RAM[16'h250B] = 8'h00;
RAM[16'h250C] = 8'h00;
RAM[16'h250D] = 8'h00;
RAM[16'h250E] = 8'h00;
RAM[16'h250F] = 8'h00;
RAM[16'h2510] = 8'h00;
RAM[16'h2511] = 8'h00;
RAM[16'h2512] = 8'h00;
RAM[16'h2513] = 8'h00;
RAM[16'h2514] = 8'h00;
RAM[16'h2515] = 8'h00;
RAM[16'h2516] = 8'h00;
RAM[16'h2517] = 8'h00;
RAM[16'h2518] = 8'h00;
RAM[16'h2519] = 8'h00;
RAM[16'h251A] = 8'h00;
RAM[16'h251B] = 8'h00;
RAM[16'h251C] = 8'h00;
RAM[16'h251D] = 8'h00;
RAM[16'h251E] = 8'h00;
RAM[16'h251F] = 8'h00;
RAM[16'h2520] = 8'h00;
RAM[16'h2521] = 8'h00;
RAM[16'h2522] = 8'h00;
RAM[16'h2523] = 8'h00;
RAM[16'h2524] = 8'h00;
RAM[16'h2525] = 8'h00;
RAM[16'h2526] = 8'h00;
RAM[16'h2527] = 8'h00;
RAM[16'h2528] = 8'h00;
RAM[16'h2529] = 8'h00;
RAM[16'h252A] = 8'h00;
RAM[16'h252B] = 8'h00;
RAM[16'h252C] = 8'h00;
RAM[16'h252D] = 8'h00;
RAM[16'h252E] = 8'h00;
RAM[16'h252F] = 8'h00;
RAM[16'h2530] = 8'h00;
RAM[16'h2531] = 8'h00;
RAM[16'h2532] = 8'h00;
RAM[16'h2533] = 8'h00;
RAM[16'h2534] = 8'h00;
RAM[16'h2535] = 8'h00;
RAM[16'h2536] = 8'h00;
RAM[16'h2537] = 8'h00;
RAM[16'h2538] = 8'h00;
RAM[16'h2539] = 8'h00;
RAM[16'h253A] = 8'h00;
RAM[16'h253B] = 8'h00;
RAM[16'h253C] = 8'h00;
RAM[16'h253D] = 8'h00;
RAM[16'h253E] = 8'h00;
RAM[16'h253F] = 8'h00;
RAM[16'h2540] = 8'h00;
RAM[16'h2541] = 8'h00;
RAM[16'h2542] = 8'h00;
RAM[16'h2543] = 8'h00;
RAM[16'h2544] = 8'h00;
RAM[16'h2545] = 8'h00;
RAM[16'h2546] = 8'h00;
RAM[16'h2547] = 8'h00;
RAM[16'h2548] = 8'h00;
RAM[16'h2549] = 8'h00;
RAM[16'h254A] = 8'h00;
RAM[16'h254B] = 8'h00;
RAM[16'h254C] = 8'h00;
RAM[16'h254D] = 8'h00;
RAM[16'h254E] = 8'h00;
RAM[16'h254F] = 8'h00;
RAM[16'h2550] = 8'h00;
RAM[16'h2551] = 8'h00;
RAM[16'h2552] = 8'h00;
RAM[16'h2553] = 8'h00;
RAM[16'h2554] = 8'h00;
RAM[16'h2555] = 8'h00;
RAM[16'h2556] = 8'h00;
RAM[16'h2557] = 8'h00;
RAM[16'h2558] = 8'h00;
RAM[16'h2559] = 8'h00;
RAM[16'h255A] = 8'h00;
RAM[16'h255B] = 8'h00;
RAM[16'h255C] = 8'h00;
RAM[16'h255D] = 8'h00;
RAM[16'h255E] = 8'h00;
RAM[16'h255F] = 8'h00;
RAM[16'h2560] = 8'h00;
RAM[16'h2561] = 8'h00;
RAM[16'h2562] = 8'h00;
RAM[16'h2563] = 8'h00;
RAM[16'h2564] = 8'h00;
RAM[16'h2565] = 8'h00;
RAM[16'h2566] = 8'h00;
RAM[16'h2567] = 8'h00;
RAM[16'h2568] = 8'h00;
RAM[16'h2569] = 8'h00;
RAM[16'h256A] = 8'h00;
RAM[16'h256B] = 8'h00;
RAM[16'h256C] = 8'h00;
RAM[16'h256D] = 8'h00;
RAM[16'h256E] = 8'h00;
RAM[16'h256F] = 8'h00;
RAM[16'h2570] = 8'h00;
RAM[16'h2571] = 8'h00;
RAM[16'h2572] = 8'h00;
RAM[16'h2573] = 8'h00;
RAM[16'h2574] = 8'h00;
RAM[16'h2575] = 8'h00;
RAM[16'h2576] = 8'h00;
RAM[16'h2577] = 8'h00;
RAM[16'h2578] = 8'h00;
RAM[16'h2579] = 8'h00;
RAM[16'h257A] = 8'h00;
RAM[16'h257B] = 8'h00;
RAM[16'h257C] = 8'h00;
RAM[16'h257D] = 8'h00;
RAM[16'h257E] = 8'h00;
RAM[16'h257F] = 8'h00;
RAM[16'h2580] = 8'h00;
RAM[16'h2581] = 8'h00;
RAM[16'h2582] = 8'h00;
RAM[16'h2583] = 8'h00;
RAM[16'h2584] = 8'h00;
RAM[16'h2585] = 8'h00;
RAM[16'h2586] = 8'h00;
RAM[16'h2587] = 8'h00;
RAM[16'h2588] = 8'h00;
RAM[16'h2589] = 8'h00;
RAM[16'h258A] = 8'h00;
RAM[16'h258B] = 8'h00;
RAM[16'h258C] = 8'h00;
RAM[16'h258D] = 8'h00;
RAM[16'h258E] = 8'h00;
RAM[16'h258F] = 8'h00;
RAM[16'h2590] = 8'h00;
RAM[16'h2591] = 8'h00;
RAM[16'h2592] = 8'h00;
RAM[16'h2593] = 8'h00;
RAM[16'h2594] = 8'h00;
RAM[16'h2595] = 8'h00;
RAM[16'h2596] = 8'h00;
RAM[16'h2597] = 8'h00;
RAM[16'h2598] = 8'h00;
RAM[16'h2599] = 8'h00;
RAM[16'h259A] = 8'h00;
RAM[16'h259B] = 8'h00;
RAM[16'h259C] = 8'h00;
RAM[16'h259D] = 8'h00;
RAM[16'h259E] = 8'h00;
RAM[16'h259F] = 8'h00;
RAM[16'h25A0] = 8'h00;
RAM[16'h25A1] = 8'h00;
RAM[16'h25A2] = 8'h00;
RAM[16'h25A3] = 8'h00;
RAM[16'h25A4] = 8'h00;
RAM[16'h25A5] = 8'h00;
RAM[16'h25A6] = 8'h00;
RAM[16'h25A7] = 8'h00;
RAM[16'h25A8] = 8'h00;
RAM[16'h25A9] = 8'h00;
RAM[16'h25AA] = 8'h00;
RAM[16'h25AB] = 8'h00;
RAM[16'h25AC] = 8'h00;
RAM[16'h25AD] = 8'h00;
RAM[16'h25AE] = 8'h00;
RAM[16'h25AF] = 8'h00;
RAM[16'h25B0] = 8'h00;
RAM[16'h25B1] = 8'h00;
RAM[16'h25B2] = 8'h00;
RAM[16'h25B3] = 8'h00;
RAM[16'h25B4] = 8'h00;
RAM[16'h25B5] = 8'h00;
RAM[16'h25B6] = 8'h00;
RAM[16'h25B7] = 8'h00;
RAM[16'h25B8] = 8'h00;
RAM[16'h25B9] = 8'h00;
RAM[16'h25BA] = 8'h00;
RAM[16'h25BB] = 8'h00;
RAM[16'h25BC] = 8'h00;
RAM[16'h25BD] = 8'h00;
RAM[16'h25BE] = 8'h00;
RAM[16'h25BF] = 8'h00;
RAM[16'h25C0] = 8'h00;
RAM[16'h25C1] = 8'h00;
RAM[16'h25C2] = 8'h00;
RAM[16'h25C3] = 8'h00;
RAM[16'h25C4] = 8'h00;
RAM[16'h25C5] = 8'h00;
RAM[16'h25C6] = 8'h00;
RAM[16'h25C7] = 8'h00;
RAM[16'h25C8] = 8'h00;
RAM[16'h25C9] = 8'h00;
RAM[16'h25CA] = 8'h00;
RAM[16'h25CB] = 8'h00;
RAM[16'h25CC] = 8'h00;
RAM[16'h25CD] = 8'h00;
RAM[16'h25CE] = 8'h00;
RAM[16'h25CF] = 8'h00;
RAM[16'h25D0] = 8'h00;
RAM[16'h25D1] = 8'h00;
RAM[16'h25D2] = 8'h00;
RAM[16'h25D3] = 8'h00;
RAM[16'h25D4] = 8'h00;
RAM[16'h25D5] = 8'h00;
RAM[16'h25D6] = 8'h00;
RAM[16'h25D7] = 8'h00;
RAM[16'h25D8] = 8'h00;
RAM[16'h25D9] = 8'h00;
RAM[16'h25DA] = 8'h00;
RAM[16'h25DB] = 8'h00;
RAM[16'h25DC] = 8'h00;
RAM[16'h25DD] = 8'h00;
RAM[16'h25DE] = 8'h00;
RAM[16'h25DF] = 8'h00;
RAM[16'h25E0] = 8'h00;
RAM[16'h25E1] = 8'h00;
RAM[16'h25E2] = 8'h00;
RAM[16'h25E3] = 8'h00;
RAM[16'h25E4] = 8'h00;
RAM[16'h25E5] = 8'h00;
RAM[16'h25E6] = 8'h00;
RAM[16'h25E7] = 8'h00;
RAM[16'h25E8] = 8'h00;
RAM[16'h25E9] = 8'h00;
RAM[16'h25EA] = 8'h00;
RAM[16'h25EB] = 8'h00;
RAM[16'h25EC] = 8'h00;
RAM[16'h25ED] = 8'h00;
RAM[16'h25EE] = 8'h00;
RAM[16'h25EF] = 8'h00;
RAM[16'h25F0] = 8'h00;
RAM[16'h25F1] = 8'h00;
RAM[16'h25F2] = 8'h00;
RAM[16'h25F3] = 8'h00;
RAM[16'h25F4] = 8'h00;
RAM[16'h25F5] = 8'h00;
RAM[16'h25F6] = 8'h00;
RAM[16'h25F7] = 8'h00;
RAM[16'h25F8] = 8'h00;
RAM[16'h25F9] = 8'h00;
RAM[16'h25FA] = 8'h00;
RAM[16'h25FB] = 8'h00;
RAM[16'h25FC] = 8'h00;
RAM[16'h25FD] = 8'h00;
RAM[16'h25FE] = 8'h00;
RAM[16'h25FF] = 8'h00;
RAM[16'h2600] = 8'h00;
RAM[16'h2601] = 8'h00;
RAM[16'h2602] = 8'h00;
RAM[16'h2603] = 8'h00;
RAM[16'h2604] = 8'h00;
RAM[16'h2605] = 8'h00;
RAM[16'h2606] = 8'h00;
RAM[16'h2607] = 8'h00;
RAM[16'h2608] = 8'h00;
RAM[16'h2609] = 8'h00;
RAM[16'h260A] = 8'h00;
RAM[16'h260B] = 8'h00;
RAM[16'h260C] = 8'h00;
RAM[16'h260D] = 8'h00;
RAM[16'h260E] = 8'h00;
RAM[16'h260F] = 8'h00;
RAM[16'h2610] = 8'h00;
RAM[16'h2611] = 8'h00;
RAM[16'h2612] = 8'h00;
RAM[16'h2613] = 8'h00;
RAM[16'h2614] = 8'h00;
RAM[16'h2615] = 8'h00;
RAM[16'h2616] = 8'h00;
RAM[16'h2617] = 8'h00;
RAM[16'h2618] = 8'h00;
RAM[16'h2619] = 8'h00;
RAM[16'h261A] = 8'h00;
RAM[16'h261B] = 8'h00;
RAM[16'h261C] = 8'h00;
RAM[16'h261D] = 8'h00;
RAM[16'h261E] = 8'h00;
RAM[16'h261F] = 8'h00;
RAM[16'h2620] = 8'h00;
RAM[16'h2621] = 8'h00;
RAM[16'h2622] = 8'h00;
RAM[16'h2623] = 8'h00;
RAM[16'h2624] = 8'h00;
RAM[16'h2625] = 8'h00;
RAM[16'h2626] = 8'h00;
RAM[16'h2627] = 8'h00;
RAM[16'h2628] = 8'h00;
RAM[16'h2629] = 8'h00;
RAM[16'h262A] = 8'h00;
RAM[16'h262B] = 8'h00;
RAM[16'h262C] = 8'h00;
RAM[16'h262D] = 8'h00;
RAM[16'h262E] = 8'h00;
RAM[16'h262F] = 8'h00;
RAM[16'h2630] = 8'h00;
RAM[16'h2631] = 8'h00;
RAM[16'h2632] = 8'h00;
RAM[16'h2633] = 8'h00;
RAM[16'h2634] = 8'h00;
RAM[16'h2635] = 8'h00;
RAM[16'h2636] = 8'h00;
RAM[16'h2637] = 8'h00;
RAM[16'h2638] = 8'h00;
RAM[16'h2639] = 8'h00;
RAM[16'h263A] = 8'h00;
RAM[16'h263B] = 8'h00;
RAM[16'h263C] = 8'h00;
RAM[16'h263D] = 8'h00;
RAM[16'h263E] = 8'h00;
RAM[16'h263F] = 8'h00;
RAM[16'h2640] = 8'h00;
RAM[16'h2641] = 8'h00;
RAM[16'h2642] = 8'h00;
RAM[16'h2643] = 8'h00;
RAM[16'h2644] = 8'h00;
RAM[16'h2645] = 8'h00;
RAM[16'h2646] = 8'h00;
RAM[16'h2647] = 8'h00;
RAM[16'h2648] = 8'h00;
RAM[16'h2649] = 8'h00;
RAM[16'h264A] = 8'h00;
RAM[16'h264B] = 8'h00;
RAM[16'h264C] = 8'h00;
RAM[16'h264D] = 8'h00;
RAM[16'h264E] = 8'h00;
RAM[16'h264F] = 8'h00;
RAM[16'h2650] = 8'h00;
RAM[16'h2651] = 8'h00;
RAM[16'h2652] = 8'h00;
RAM[16'h2653] = 8'h00;
RAM[16'h2654] = 8'h00;
RAM[16'h2655] = 8'h00;
RAM[16'h2656] = 8'h00;
RAM[16'h2657] = 8'h00;
RAM[16'h2658] = 8'h00;
RAM[16'h2659] = 8'h00;
RAM[16'h265A] = 8'h00;
RAM[16'h265B] = 8'h00;
RAM[16'h265C] = 8'h00;
RAM[16'h265D] = 8'h00;
RAM[16'h265E] = 8'h00;
RAM[16'h265F] = 8'h00;
RAM[16'h2660] = 8'h00;
RAM[16'h2661] = 8'h00;
RAM[16'h2662] = 8'h00;
RAM[16'h2663] = 8'h00;
RAM[16'h2664] = 8'h00;
RAM[16'h2665] = 8'h00;
RAM[16'h2666] = 8'h00;
RAM[16'h2667] = 8'h00;
RAM[16'h2668] = 8'h00;
RAM[16'h2669] = 8'h00;
RAM[16'h266A] = 8'h00;
RAM[16'h266B] = 8'h00;
RAM[16'h266C] = 8'h00;
RAM[16'h266D] = 8'h00;
RAM[16'h266E] = 8'h00;
RAM[16'h266F] = 8'h00;
RAM[16'h2670] = 8'h00;
RAM[16'h2671] = 8'h00;
RAM[16'h2672] = 8'h00;
RAM[16'h2673] = 8'h00;
RAM[16'h2674] = 8'h00;
RAM[16'h2675] = 8'h00;
RAM[16'h2676] = 8'h00;
RAM[16'h2677] = 8'h00;
RAM[16'h2678] = 8'h00;
RAM[16'h2679] = 8'h00;
RAM[16'h267A] = 8'h00;
RAM[16'h267B] = 8'h00;
RAM[16'h267C] = 8'h00;
RAM[16'h267D] = 8'h00;
RAM[16'h267E] = 8'h00;
RAM[16'h267F] = 8'h00;
RAM[16'h2680] = 8'h00;
RAM[16'h2681] = 8'h00;
RAM[16'h2682] = 8'h00;
RAM[16'h2683] = 8'h00;
RAM[16'h2684] = 8'h00;
RAM[16'h2685] = 8'h00;
RAM[16'h2686] = 8'h00;
RAM[16'h2687] = 8'h00;
RAM[16'h2688] = 8'h00;
RAM[16'h2689] = 8'h00;
RAM[16'h268A] = 8'h00;
RAM[16'h268B] = 8'h00;
RAM[16'h268C] = 8'h00;
RAM[16'h268D] = 8'h00;
RAM[16'h268E] = 8'h00;
RAM[16'h268F] = 8'h00;
RAM[16'h2690] = 8'h00;
RAM[16'h2691] = 8'h00;
RAM[16'h2692] = 8'h00;
RAM[16'h2693] = 8'h00;
RAM[16'h2694] = 8'h00;
RAM[16'h2695] = 8'h00;
RAM[16'h2696] = 8'h00;
RAM[16'h2697] = 8'h00;
RAM[16'h2698] = 8'h00;
RAM[16'h2699] = 8'h00;
RAM[16'h269A] = 8'h00;
RAM[16'h269B] = 8'h00;
RAM[16'h269C] = 8'h00;
RAM[16'h269D] = 8'h00;
RAM[16'h269E] = 8'h00;
RAM[16'h269F] = 8'h00;
RAM[16'h26A0] = 8'h00;
RAM[16'h26A1] = 8'h00;
RAM[16'h26A2] = 8'h00;
RAM[16'h26A3] = 8'h00;
RAM[16'h26A4] = 8'h00;
RAM[16'h26A5] = 8'h00;
RAM[16'h26A6] = 8'h00;
RAM[16'h26A7] = 8'h00;
RAM[16'h26A8] = 8'h00;
RAM[16'h26A9] = 8'h00;
RAM[16'h26AA] = 8'h00;
RAM[16'h26AB] = 8'h00;
RAM[16'h26AC] = 8'h00;
RAM[16'h26AD] = 8'h00;
RAM[16'h26AE] = 8'h00;
RAM[16'h26AF] = 8'h00;
RAM[16'h26B0] = 8'h00;
RAM[16'h26B1] = 8'h00;
RAM[16'h26B2] = 8'h00;
RAM[16'h26B3] = 8'h00;
RAM[16'h26B4] = 8'h00;
RAM[16'h26B5] = 8'h00;
RAM[16'h26B6] = 8'h00;
RAM[16'h26B7] = 8'h00;
RAM[16'h26B8] = 8'h00;
RAM[16'h26B9] = 8'h00;
RAM[16'h26BA] = 8'h00;
RAM[16'h26BB] = 8'h00;
RAM[16'h26BC] = 8'h00;
RAM[16'h26BD] = 8'h00;
RAM[16'h26BE] = 8'h00;
RAM[16'h26BF] = 8'h00;
RAM[16'h26C0] = 8'h00;
RAM[16'h26C1] = 8'h00;
RAM[16'h26C2] = 8'h00;
RAM[16'h26C3] = 8'h00;
RAM[16'h26C4] = 8'h00;
RAM[16'h26C5] = 8'h00;
RAM[16'h26C6] = 8'h00;
RAM[16'h26C7] = 8'h00;
RAM[16'h26C8] = 8'h00;
RAM[16'h26C9] = 8'h00;
RAM[16'h26CA] = 8'h00;
RAM[16'h26CB] = 8'h00;
RAM[16'h26CC] = 8'h00;
RAM[16'h26CD] = 8'h00;
RAM[16'h26CE] = 8'h00;
RAM[16'h26CF] = 8'h00;
RAM[16'h26D0] = 8'h00;
RAM[16'h26D1] = 8'h00;
RAM[16'h26D2] = 8'h00;
RAM[16'h26D3] = 8'h00;
RAM[16'h26D4] = 8'h00;
RAM[16'h26D5] = 8'h00;
RAM[16'h26D6] = 8'h00;
RAM[16'h26D7] = 8'h00;
RAM[16'h26D8] = 8'h00;
RAM[16'h26D9] = 8'h00;
RAM[16'h26DA] = 8'h00;
RAM[16'h26DB] = 8'h00;
RAM[16'h26DC] = 8'h00;
RAM[16'h26DD] = 8'h00;
RAM[16'h26DE] = 8'h00;
RAM[16'h26DF] = 8'h00;
RAM[16'h26E0] = 8'h00;
RAM[16'h26E1] = 8'h00;
RAM[16'h26E2] = 8'h00;
RAM[16'h26E3] = 8'h00;
RAM[16'h26E4] = 8'h00;
RAM[16'h26E5] = 8'h00;
RAM[16'h26E6] = 8'h00;
RAM[16'h26E7] = 8'h00;
RAM[16'h26E8] = 8'h00;
RAM[16'h26E9] = 8'h00;
RAM[16'h26EA] = 8'h00;
RAM[16'h26EB] = 8'h00;
RAM[16'h26EC] = 8'h00;
RAM[16'h26ED] = 8'h00;
RAM[16'h26EE] = 8'h00;
RAM[16'h26EF] = 8'h00;
RAM[16'h26F0] = 8'h00;
RAM[16'h26F1] = 8'h00;
RAM[16'h26F2] = 8'h00;
RAM[16'h26F3] = 8'h00;
RAM[16'h26F4] = 8'h00;
RAM[16'h26F5] = 8'h00;
RAM[16'h26F6] = 8'h00;
RAM[16'h26F7] = 8'h00;
RAM[16'h26F8] = 8'h00;
RAM[16'h26F9] = 8'h00;
RAM[16'h26FA] = 8'h00;
RAM[16'h26FB] = 8'h00;
RAM[16'h26FC] = 8'h00;
RAM[16'h26FD] = 8'h00;
RAM[16'h26FE] = 8'h00;
RAM[16'h26FF] = 8'h00;
RAM[16'h2700] = 8'h00;
RAM[16'h2701] = 8'h00;
RAM[16'h2702] = 8'h00;
RAM[16'h2703] = 8'h00;
RAM[16'h2704] = 8'h00;
RAM[16'h2705] = 8'h00;
RAM[16'h2706] = 8'h00;
RAM[16'h2707] = 8'h00;
RAM[16'h2708] = 8'h00;
RAM[16'h2709] = 8'h00;
RAM[16'h270A] = 8'h00;
RAM[16'h270B] = 8'h00;
RAM[16'h270C] = 8'h00;
RAM[16'h270D] = 8'h00;
RAM[16'h270E] = 8'h00;
RAM[16'h270F] = 8'h00;
RAM[16'h2710] = 8'h00;
RAM[16'h2711] = 8'h00;
RAM[16'h2712] = 8'h00;
RAM[16'h2713] = 8'h00;
RAM[16'h2714] = 8'h00;
RAM[16'h2715] = 8'h00;
RAM[16'h2716] = 8'h00;
RAM[16'h2717] = 8'h00;
RAM[16'h2718] = 8'h00;
RAM[16'h2719] = 8'h00;
RAM[16'h271A] = 8'h00;
RAM[16'h271B] = 8'h00;
RAM[16'h271C] = 8'h00;
RAM[16'h271D] = 8'h00;
RAM[16'h271E] = 8'h00;
RAM[16'h271F] = 8'h00;
RAM[16'h2720] = 8'h00;
RAM[16'h2721] = 8'h00;
RAM[16'h2722] = 8'h00;
RAM[16'h2723] = 8'h00;
RAM[16'h2724] = 8'h00;
RAM[16'h2725] = 8'h00;
RAM[16'h2726] = 8'h00;
RAM[16'h2727] = 8'h00;
RAM[16'h2728] = 8'h00;
RAM[16'h2729] = 8'h00;
RAM[16'h272A] = 8'h00;
RAM[16'h272B] = 8'h00;
RAM[16'h272C] = 8'h00;
RAM[16'h272D] = 8'h00;
RAM[16'h272E] = 8'h00;
RAM[16'h272F] = 8'h00;
RAM[16'h2730] = 8'h00;
RAM[16'h2731] = 8'h00;
RAM[16'h2732] = 8'h00;
RAM[16'h2733] = 8'h00;
RAM[16'h2734] = 8'h00;
RAM[16'h2735] = 8'h00;
RAM[16'h2736] = 8'h00;
RAM[16'h2737] = 8'h00;
RAM[16'h2738] = 8'h00;
RAM[16'h2739] = 8'h00;
RAM[16'h273A] = 8'h00;
RAM[16'h273B] = 8'h00;
RAM[16'h273C] = 8'h00;
RAM[16'h273D] = 8'h00;
RAM[16'h273E] = 8'h00;
RAM[16'h273F] = 8'h00;
RAM[16'h2740] = 8'h00;
RAM[16'h2741] = 8'h00;
RAM[16'h2742] = 8'h00;
RAM[16'h2743] = 8'h00;
RAM[16'h2744] = 8'h00;
RAM[16'h2745] = 8'h00;
RAM[16'h2746] = 8'h00;
RAM[16'h2747] = 8'h00;
RAM[16'h2748] = 8'h00;
RAM[16'h2749] = 8'h00;
RAM[16'h274A] = 8'h00;
RAM[16'h274B] = 8'h00;
RAM[16'h274C] = 8'h00;
RAM[16'h274D] = 8'h00;
RAM[16'h274E] = 8'h00;
RAM[16'h274F] = 8'h00;
RAM[16'h2750] = 8'h00;
RAM[16'h2751] = 8'h00;
RAM[16'h2752] = 8'h00;
RAM[16'h2753] = 8'h00;
RAM[16'h2754] = 8'h00;
RAM[16'h2755] = 8'h00;
RAM[16'h2756] = 8'h00;
RAM[16'h2757] = 8'h00;
RAM[16'h2758] = 8'h00;
RAM[16'h2759] = 8'h00;
RAM[16'h275A] = 8'h00;
RAM[16'h275B] = 8'h00;
RAM[16'h275C] = 8'h00;
RAM[16'h275D] = 8'h00;
RAM[16'h275E] = 8'h00;
RAM[16'h275F] = 8'h00;
RAM[16'h2760] = 8'h00;
RAM[16'h2761] = 8'h00;
RAM[16'h2762] = 8'h00;
RAM[16'h2763] = 8'h00;
RAM[16'h2764] = 8'h00;
RAM[16'h2765] = 8'h00;
RAM[16'h2766] = 8'h00;
RAM[16'h2767] = 8'h00;
RAM[16'h2768] = 8'h00;
RAM[16'h2769] = 8'h00;
RAM[16'h276A] = 8'h00;
RAM[16'h276B] = 8'h00;
RAM[16'h276C] = 8'h00;
RAM[16'h276D] = 8'h00;
RAM[16'h276E] = 8'h00;
RAM[16'h276F] = 8'h00;
RAM[16'h2770] = 8'h00;
RAM[16'h2771] = 8'h00;
RAM[16'h2772] = 8'h00;
RAM[16'h2773] = 8'h00;
RAM[16'h2774] = 8'h00;
RAM[16'h2775] = 8'h00;
RAM[16'h2776] = 8'h00;
RAM[16'h2777] = 8'h00;
RAM[16'h2778] = 8'h00;
RAM[16'h2779] = 8'h00;
RAM[16'h277A] = 8'h00;
RAM[16'h277B] = 8'h00;
RAM[16'h277C] = 8'h00;
RAM[16'h277D] = 8'h00;
RAM[16'h277E] = 8'h00;
RAM[16'h277F] = 8'h00;
RAM[16'h2780] = 8'h00;
RAM[16'h2781] = 8'h00;
RAM[16'h2782] = 8'h00;
RAM[16'h2783] = 8'h00;
RAM[16'h2784] = 8'h00;
RAM[16'h2785] = 8'h00;
RAM[16'h2786] = 8'h00;
RAM[16'h2787] = 8'h00;
RAM[16'h2788] = 8'h00;
RAM[16'h2789] = 8'h00;
RAM[16'h278A] = 8'h00;
RAM[16'h278B] = 8'h00;
RAM[16'h278C] = 8'h00;
RAM[16'h278D] = 8'h00;
RAM[16'h278E] = 8'h00;
RAM[16'h278F] = 8'h00;
RAM[16'h2790] = 8'h00;
RAM[16'h2791] = 8'h00;
RAM[16'h2792] = 8'h00;
RAM[16'h2793] = 8'h00;
RAM[16'h2794] = 8'h00;
RAM[16'h2795] = 8'h00;
RAM[16'h2796] = 8'h00;
RAM[16'h2797] = 8'h00;
RAM[16'h2798] = 8'h00;
RAM[16'h2799] = 8'h00;
RAM[16'h279A] = 8'h00;
RAM[16'h279B] = 8'h00;
RAM[16'h279C] = 8'h00;
RAM[16'h279D] = 8'h00;
RAM[16'h279E] = 8'h00;
RAM[16'h279F] = 8'h00;
RAM[16'h27A0] = 8'h00;
RAM[16'h27A1] = 8'h00;
RAM[16'h27A2] = 8'h00;
RAM[16'h27A3] = 8'h00;
RAM[16'h27A4] = 8'h00;
RAM[16'h27A5] = 8'h00;
RAM[16'h27A6] = 8'h00;
RAM[16'h27A7] = 8'h00;
RAM[16'h27A8] = 8'h00;
RAM[16'h27A9] = 8'h00;
RAM[16'h27AA] = 8'h00;
RAM[16'h27AB] = 8'h00;
RAM[16'h27AC] = 8'h00;
RAM[16'h27AD] = 8'h00;
RAM[16'h27AE] = 8'h00;
RAM[16'h27AF] = 8'h00;
RAM[16'h27B0] = 8'h00;
RAM[16'h27B1] = 8'h00;
RAM[16'h27B2] = 8'h00;
RAM[16'h27B3] = 8'h00;
RAM[16'h27B4] = 8'h00;
RAM[16'h27B5] = 8'h00;
RAM[16'h27B6] = 8'h00;
RAM[16'h27B7] = 8'h00;
RAM[16'h27B8] = 8'h00;
RAM[16'h27B9] = 8'h00;
RAM[16'h27BA] = 8'h00;
RAM[16'h27BB] = 8'h00;
RAM[16'h27BC] = 8'h00;
RAM[16'h27BD] = 8'h00;
RAM[16'h27BE] = 8'h00;
RAM[16'h27BF] = 8'h00;
RAM[16'h27C0] = 8'h00;
RAM[16'h27C1] = 8'h00;
RAM[16'h27C2] = 8'h00;
RAM[16'h27C3] = 8'h00;
RAM[16'h27C4] = 8'h00;
RAM[16'h27C5] = 8'h00;
RAM[16'h27C6] = 8'h00;
RAM[16'h27C7] = 8'h00;
RAM[16'h27C8] = 8'h00;
RAM[16'h27C9] = 8'h00;
RAM[16'h27CA] = 8'h00;
RAM[16'h27CB] = 8'h00;
RAM[16'h27CC] = 8'h00;
RAM[16'h27CD] = 8'h00;
RAM[16'h27CE] = 8'h00;
RAM[16'h27CF] = 8'h00;
RAM[16'h27D0] = 8'h00;
RAM[16'h27D1] = 8'h00;
RAM[16'h27D2] = 8'h00;
RAM[16'h27D3] = 8'h00;
RAM[16'h27D4] = 8'h00;
RAM[16'h27D5] = 8'h00;
RAM[16'h27D6] = 8'h00;
RAM[16'h27D7] = 8'h00;
RAM[16'h27D8] = 8'h00;
RAM[16'h27D9] = 8'h00;
RAM[16'h27DA] = 8'h00;
RAM[16'h27DB] = 8'h00;
RAM[16'h27DC] = 8'h00;
RAM[16'h27DD] = 8'h00;
RAM[16'h27DE] = 8'h00;
RAM[16'h27DF] = 8'h00;
RAM[16'h27E0] = 8'h00;
RAM[16'h27E1] = 8'h00;
RAM[16'h27E2] = 8'h00;
RAM[16'h27E3] = 8'h00;
RAM[16'h27E4] = 8'h00;
RAM[16'h27E5] = 8'h00;
RAM[16'h27E6] = 8'h00;
RAM[16'h27E7] = 8'h00;
RAM[16'h27E8] = 8'h00;
RAM[16'h27E9] = 8'h00;
RAM[16'h27EA] = 8'h00;
RAM[16'h27EB] = 8'h00;
RAM[16'h27EC] = 8'h00;
RAM[16'h27ED] = 8'h00;
RAM[16'h27EE] = 8'h00;
RAM[16'h27EF] = 8'h00;
RAM[16'h27F0] = 8'h00;
RAM[16'h27F1] = 8'h00;
RAM[16'h27F2] = 8'h00;
RAM[16'h27F3] = 8'h00;
RAM[16'h27F4] = 8'h00;
RAM[16'h27F5] = 8'h00;
RAM[16'h27F6] = 8'h00;
RAM[16'h27F7] = 8'h00;
RAM[16'h27F8] = 8'h00;
RAM[16'h27F9] = 8'h00;
RAM[16'h27FA] = 8'h00;
RAM[16'h27FB] = 8'h00;
RAM[16'h27FC] = 8'h00;
RAM[16'h27FD] = 8'h00;
RAM[16'h27FE] = 8'h00;
RAM[16'h27FF] = 8'h00;
RAM[16'h2800] = 8'h00;
RAM[16'h2801] = 8'h00;
RAM[16'h2802] = 8'h00;
RAM[16'h2803] = 8'h00;
RAM[16'h2804] = 8'h00;
RAM[16'h2805] = 8'h00;
RAM[16'h2806] = 8'h00;
RAM[16'h2807] = 8'h00;
RAM[16'h2808] = 8'h00;
RAM[16'h2809] = 8'h00;
RAM[16'h280A] = 8'h00;
RAM[16'h280B] = 8'h00;
RAM[16'h280C] = 8'h00;
RAM[16'h280D] = 8'h00;
RAM[16'h280E] = 8'h00;
RAM[16'h280F] = 8'h00;
RAM[16'h2810] = 8'h00;
RAM[16'h2811] = 8'h00;
RAM[16'h2812] = 8'h00;
RAM[16'h2813] = 8'h00;
RAM[16'h2814] = 8'h00;
RAM[16'h2815] = 8'h00;
RAM[16'h2816] = 8'h00;
RAM[16'h2817] = 8'h00;
RAM[16'h2818] = 8'h00;
RAM[16'h2819] = 8'h00;
RAM[16'h281A] = 8'h00;
RAM[16'h281B] = 8'h00;
RAM[16'h281C] = 8'h00;
RAM[16'h281D] = 8'h00;
RAM[16'h281E] = 8'h00;
RAM[16'h281F] = 8'h00;
RAM[16'h2820] = 8'h00;
RAM[16'h2821] = 8'h00;
RAM[16'h2822] = 8'h00;
RAM[16'h2823] = 8'h00;
RAM[16'h2824] = 8'h00;
RAM[16'h2825] = 8'h00;
RAM[16'h2826] = 8'h00;
RAM[16'h2827] = 8'h00;
RAM[16'h2828] = 8'h00;
RAM[16'h2829] = 8'h00;
RAM[16'h282A] = 8'h00;
RAM[16'h282B] = 8'h00;
RAM[16'h282C] = 8'h00;
RAM[16'h282D] = 8'h00;
RAM[16'h282E] = 8'h00;
RAM[16'h282F] = 8'h00;
RAM[16'h2830] = 8'h00;
RAM[16'h2831] = 8'h00;
RAM[16'h2832] = 8'h00;
RAM[16'h2833] = 8'h00;
RAM[16'h2834] = 8'h00;
RAM[16'h2835] = 8'h00;
RAM[16'h2836] = 8'h00;
RAM[16'h2837] = 8'h00;
RAM[16'h2838] = 8'h00;
RAM[16'h2839] = 8'h00;
RAM[16'h283A] = 8'h00;
RAM[16'h283B] = 8'h00;
RAM[16'h283C] = 8'h00;
RAM[16'h283D] = 8'h00;
RAM[16'h283E] = 8'h00;
RAM[16'h283F] = 8'h00;
RAM[16'h2840] = 8'h00;
RAM[16'h2841] = 8'h00;
RAM[16'h2842] = 8'h00;
RAM[16'h2843] = 8'h00;
RAM[16'h2844] = 8'h00;
RAM[16'h2845] = 8'h00;
RAM[16'h2846] = 8'h00;
RAM[16'h2847] = 8'h00;
RAM[16'h2848] = 8'h00;
RAM[16'h2849] = 8'h00;
RAM[16'h284A] = 8'h00;
RAM[16'h284B] = 8'h00;
RAM[16'h284C] = 8'h00;
RAM[16'h284D] = 8'h00;
RAM[16'h284E] = 8'h00;
RAM[16'h284F] = 8'h00;
RAM[16'h2850] = 8'h00;
RAM[16'h2851] = 8'h00;
RAM[16'h2852] = 8'h00;
RAM[16'h2853] = 8'h00;
RAM[16'h2854] = 8'h00;
RAM[16'h2855] = 8'h00;
RAM[16'h2856] = 8'h00;
RAM[16'h2857] = 8'h00;
RAM[16'h2858] = 8'h00;
RAM[16'h2859] = 8'h00;
RAM[16'h285A] = 8'h00;
RAM[16'h285B] = 8'h00;
RAM[16'h285C] = 8'h00;
RAM[16'h285D] = 8'h00;
RAM[16'h285E] = 8'h00;
RAM[16'h285F] = 8'h00;
RAM[16'h2860] = 8'h00;
RAM[16'h2861] = 8'h00;
RAM[16'h2862] = 8'h00;
RAM[16'h2863] = 8'h00;
RAM[16'h2864] = 8'h00;
RAM[16'h2865] = 8'h00;
RAM[16'h2866] = 8'h00;
RAM[16'h2867] = 8'h00;
RAM[16'h2868] = 8'h00;
RAM[16'h2869] = 8'h00;
RAM[16'h286A] = 8'h00;
RAM[16'h286B] = 8'h00;
RAM[16'h286C] = 8'h00;
RAM[16'h286D] = 8'h00;
RAM[16'h286E] = 8'h00;
RAM[16'h286F] = 8'h00;
RAM[16'h2870] = 8'h00;
RAM[16'h2871] = 8'h00;
RAM[16'h2872] = 8'h00;
RAM[16'h2873] = 8'h00;
RAM[16'h2874] = 8'h00;
RAM[16'h2875] = 8'h00;
RAM[16'h2876] = 8'h00;
RAM[16'h2877] = 8'h00;
RAM[16'h2878] = 8'h00;
RAM[16'h2879] = 8'h00;
RAM[16'h287A] = 8'h00;
RAM[16'h287B] = 8'h00;
RAM[16'h287C] = 8'h00;
RAM[16'h287D] = 8'h00;
RAM[16'h287E] = 8'h00;
RAM[16'h287F] = 8'h00;
RAM[16'h2880] = 8'h00;
RAM[16'h2881] = 8'h00;
RAM[16'h2882] = 8'h00;
RAM[16'h2883] = 8'h00;
RAM[16'h2884] = 8'h00;
RAM[16'h2885] = 8'h00;
RAM[16'h2886] = 8'h00;
RAM[16'h2887] = 8'h00;
RAM[16'h2888] = 8'h00;
RAM[16'h2889] = 8'h00;
RAM[16'h288A] = 8'h00;
RAM[16'h288B] = 8'h00;
RAM[16'h288C] = 8'h00;
RAM[16'h288D] = 8'h00;
RAM[16'h288E] = 8'h00;
RAM[16'h288F] = 8'h00;
RAM[16'h2890] = 8'h00;
RAM[16'h2891] = 8'h00;
RAM[16'h2892] = 8'h00;
RAM[16'h2893] = 8'h00;
RAM[16'h2894] = 8'h00;
RAM[16'h2895] = 8'h00;
RAM[16'h2896] = 8'h00;
RAM[16'h2897] = 8'h00;
RAM[16'h2898] = 8'h00;
RAM[16'h2899] = 8'h00;
RAM[16'h289A] = 8'h00;
RAM[16'h289B] = 8'h00;
RAM[16'h289C] = 8'h00;
RAM[16'h289D] = 8'h00;
RAM[16'h289E] = 8'h00;
RAM[16'h289F] = 8'h00;
RAM[16'h28A0] = 8'h00;
RAM[16'h28A1] = 8'h00;
RAM[16'h28A2] = 8'h00;
RAM[16'h28A3] = 8'h00;
RAM[16'h28A4] = 8'h00;
RAM[16'h28A5] = 8'h00;
RAM[16'h28A6] = 8'h00;
RAM[16'h28A7] = 8'h00;
RAM[16'h28A8] = 8'h00;
RAM[16'h28A9] = 8'h00;
RAM[16'h28AA] = 8'h00;
RAM[16'h28AB] = 8'h00;
RAM[16'h28AC] = 8'h00;
RAM[16'h28AD] = 8'h00;
RAM[16'h28AE] = 8'h00;
RAM[16'h28AF] = 8'h00;
RAM[16'h28B0] = 8'h00;
RAM[16'h28B1] = 8'h00;
RAM[16'h28B2] = 8'h00;
RAM[16'h28B3] = 8'h00;
RAM[16'h28B4] = 8'h00;
RAM[16'h28B5] = 8'h00;
RAM[16'h28B6] = 8'h00;
RAM[16'h28B7] = 8'h00;
RAM[16'h28B8] = 8'h00;
RAM[16'h28B9] = 8'h00;
RAM[16'h28BA] = 8'h00;
RAM[16'h28BB] = 8'h00;
RAM[16'h28BC] = 8'h00;
RAM[16'h28BD] = 8'h00;
RAM[16'h28BE] = 8'h00;
RAM[16'h28BF] = 8'h00;
RAM[16'h28C0] = 8'h00;
RAM[16'h28C1] = 8'h00;
RAM[16'h28C2] = 8'h00;
RAM[16'h28C3] = 8'h00;
RAM[16'h28C4] = 8'h00;
RAM[16'h28C5] = 8'h00;
RAM[16'h28C6] = 8'h00;
RAM[16'h28C7] = 8'h00;
RAM[16'h28C8] = 8'h00;
RAM[16'h28C9] = 8'h00;
RAM[16'h28CA] = 8'h00;
RAM[16'h28CB] = 8'h00;
RAM[16'h28CC] = 8'h00;
RAM[16'h28CD] = 8'h00;
RAM[16'h28CE] = 8'h00;
RAM[16'h28CF] = 8'h00;
RAM[16'h28D0] = 8'h00;
RAM[16'h28D1] = 8'h00;
RAM[16'h28D2] = 8'h00;
RAM[16'h28D3] = 8'h00;
RAM[16'h28D4] = 8'h00;
RAM[16'h28D5] = 8'h00;
RAM[16'h28D6] = 8'h00;
RAM[16'h28D7] = 8'h00;
RAM[16'h28D8] = 8'h00;
RAM[16'h28D9] = 8'h00;
RAM[16'h28DA] = 8'h00;
RAM[16'h28DB] = 8'h00;
RAM[16'h28DC] = 8'h00;
RAM[16'h28DD] = 8'h00;
RAM[16'h28DE] = 8'h00;
RAM[16'h28DF] = 8'h00;
RAM[16'h28E0] = 8'h00;
RAM[16'h28E1] = 8'h00;
RAM[16'h28E2] = 8'h00;
RAM[16'h28E3] = 8'h00;
RAM[16'h28E4] = 8'h00;
RAM[16'h28E5] = 8'h00;
RAM[16'h28E6] = 8'h00;
RAM[16'h28E7] = 8'h00;
RAM[16'h28E8] = 8'h00;
RAM[16'h28E9] = 8'h00;
RAM[16'h28EA] = 8'h00;
RAM[16'h28EB] = 8'h00;
RAM[16'h28EC] = 8'h00;
RAM[16'h28ED] = 8'h00;
RAM[16'h28EE] = 8'h00;
RAM[16'h28EF] = 8'h00;
RAM[16'h28F0] = 8'h00;
RAM[16'h28F1] = 8'h00;
RAM[16'h28F2] = 8'h00;
RAM[16'h28F3] = 8'h00;
RAM[16'h28F4] = 8'h00;
RAM[16'h28F5] = 8'h00;
RAM[16'h28F6] = 8'h00;
RAM[16'h28F7] = 8'h00;
RAM[16'h28F8] = 8'h00;
RAM[16'h28F9] = 8'h00;
RAM[16'h28FA] = 8'h00;
RAM[16'h28FB] = 8'h00;
RAM[16'h28FC] = 8'h00;
RAM[16'h28FD] = 8'h00;
RAM[16'h28FE] = 8'h00;
RAM[16'h28FF] = 8'h00;
RAM[16'h2900] = 8'h00;
RAM[16'h2901] = 8'h00;
RAM[16'h2902] = 8'h00;
RAM[16'h2903] = 8'h00;
RAM[16'h2904] = 8'h00;
RAM[16'h2905] = 8'h00;
RAM[16'h2906] = 8'h00;
RAM[16'h2907] = 8'h00;
RAM[16'h2908] = 8'h00;
RAM[16'h2909] = 8'h00;
RAM[16'h290A] = 8'h00;
RAM[16'h290B] = 8'h00;
RAM[16'h290C] = 8'h00;
RAM[16'h290D] = 8'h00;
RAM[16'h290E] = 8'h00;
RAM[16'h290F] = 8'h00;
RAM[16'h2910] = 8'h00;
RAM[16'h2911] = 8'h00;
RAM[16'h2912] = 8'h00;
RAM[16'h2913] = 8'h00;
RAM[16'h2914] = 8'h00;
RAM[16'h2915] = 8'h00;
RAM[16'h2916] = 8'h00;
RAM[16'h2917] = 8'h00;
RAM[16'h2918] = 8'h00;
RAM[16'h2919] = 8'h00;
RAM[16'h291A] = 8'h00;
RAM[16'h291B] = 8'h00;
RAM[16'h291C] = 8'h00;
RAM[16'h291D] = 8'h00;
RAM[16'h291E] = 8'h00;
RAM[16'h291F] = 8'h00;
RAM[16'h2920] = 8'h00;
RAM[16'h2921] = 8'h00;
RAM[16'h2922] = 8'h00;
RAM[16'h2923] = 8'h00;
RAM[16'h2924] = 8'h00;
RAM[16'h2925] = 8'h00;
RAM[16'h2926] = 8'h00;
RAM[16'h2927] = 8'h00;
RAM[16'h2928] = 8'h00;
RAM[16'h2929] = 8'h00;
RAM[16'h292A] = 8'h00;
RAM[16'h292B] = 8'h00;
RAM[16'h292C] = 8'h00;
RAM[16'h292D] = 8'h00;
RAM[16'h292E] = 8'h00;
RAM[16'h292F] = 8'h00;
RAM[16'h2930] = 8'h00;
RAM[16'h2931] = 8'h00;
RAM[16'h2932] = 8'h00;
RAM[16'h2933] = 8'h00;
RAM[16'h2934] = 8'h00;
RAM[16'h2935] = 8'h00;
RAM[16'h2936] = 8'h00;
RAM[16'h2937] = 8'h00;
RAM[16'h2938] = 8'h00;
RAM[16'h2939] = 8'h00;
RAM[16'h293A] = 8'h00;
RAM[16'h293B] = 8'h00;
RAM[16'h293C] = 8'h00;
RAM[16'h293D] = 8'h00;
RAM[16'h293E] = 8'h00;
RAM[16'h293F] = 8'h00;
RAM[16'h2940] = 8'h00;
RAM[16'h2941] = 8'h00;
RAM[16'h2942] = 8'h00;
RAM[16'h2943] = 8'h00;
RAM[16'h2944] = 8'h00;
RAM[16'h2945] = 8'h00;
RAM[16'h2946] = 8'h00;
RAM[16'h2947] = 8'h00;
RAM[16'h2948] = 8'h00;
RAM[16'h2949] = 8'h00;
RAM[16'h294A] = 8'h00;
RAM[16'h294B] = 8'h00;
RAM[16'h294C] = 8'h00;
RAM[16'h294D] = 8'h00;
RAM[16'h294E] = 8'h00;
RAM[16'h294F] = 8'h00;
RAM[16'h2950] = 8'h00;
RAM[16'h2951] = 8'h00;
RAM[16'h2952] = 8'h00;
RAM[16'h2953] = 8'h00;
RAM[16'h2954] = 8'h00;
RAM[16'h2955] = 8'h00;
RAM[16'h2956] = 8'h00;
RAM[16'h2957] = 8'h00;
RAM[16'h2958] = 8'h00;
RAM[16'h2959] = 8'h00;
RAM[16'h295A] = 8'h00;
RAM[16'h295B] = 8'h00;
RAM[16'h295C] = 8'h00;
RAM[16'h295D] = 8'h00;
RAM[16'h295E] = 8'h00;
RAM[16'h295F] = 8'h00;
RAM[16'h2960] = 8'h00;
RAM[16'h2961] = 8'h00;
RAM[16'h2962] = 8'h00;
RAM[16'h2963] = 8'h00;
RAM[16'h2964] = 8'h00;
RAM[16'h2965] = 8'h00;
RAM[16'h2966] = 8'h00;
RAM[16'h2967] = 8'h00;
RAM[16'h2968] = 8'h00;
RAM[16'h2969] = 8'h00;
RAM[16'h296A] = 8'h00;
RAM[16'h296B] = 8'h00;
RAM[16'h296C] = 8'h00;
RAM[16'h296D] = 8'h00;
RAM[16'h296E] = 8'h00;
RAM[16'h296F] = 8'h00;
RAM[16'h2970] = 8'h00;
RAM[16'h2971] = 8'h00;
RAM[16'h2972] = 8'h00;
RAM[16'h2973] = 8'h00;
RAM[16'h2974] = 8'h00;
RAM[16'h2975] = 8'h00;
RAM[16'h2976] = 8'h00;
RAM[16'h2977] = 8'h00;
RAM[16'h2978] = 8'h00;
RAM[16'h2979] = 8'h00;
RAM[16'h297A] = 8'h00;
RAM[16'h297B] = 8'h00;
RAM[16'h297C] = 8'h00;
RAM[16'h297D] = 8'h00;
RAM[16'h297E] = 8'h00;
RAM[16'h297F] = 8'h00;
RAM[16'h2980] = 8'h00;
RAM[16'h2981] = 8'h00;
RAM[16'h2982] = 8'h00;
RAM[16'h2983] = 8'h00;
RAM[16'h2984] = 8'h00;
RAM[16'h2985] = 8'h00;
RAM[16'h2986] = 8'h00;
RAM[16'h2987] = 8'h00;
RAM[16'h2988] = 8'h00;
RAM[16'h2989] = 8'h00;
RAM[16'h298A] = 8'h00;
RAM[16'h298B] = 8'h00;
RAM[16'h298C] = 8'h00;
RAM[16'h298D] = 8'h00;
RAM[16'h298E] = 8'h00;
RAM[16'h298F] = 8'h00;
RAM[16'h2990] = 8'h00;
RAM[16'h2991] = 8'h00;
RAM[16'h2992] = 8'h00;
RAM[16'h2993] = 8'h00;
RAM[16'h2994] = 8'h00;
RAM[16'h2995] = 8'h00;
RAM[16'h2996] = 8'h00;
RAM[16'h2997] = 8'h00;
RAM[16'h2998] = 8'h00;
RAM[16'h2999] = 8'h00;
RAM[16'h299A] = 8'h00;
RAM[16'h299B] = 8'h00;
RAM[16'h299C] = 8'h00;
RAM[16'h299D] = 8'h00;
RAM[16'h299E] = 8'h00;
RAM[16'h299F] = 8'h00;
RAM[16'h29A0] = 8'h00;
RAM[16'h29A1] = 8'h00;
RAM[16'h29A2] = 8'h00;
RAM[16'h29A3] = 8'h00;
RAM[16'h29A4] = 8'h00;
RAM[16'h29A5] = 8'h00;
RAM[16'h29A6] = 8'h00;
RAM[16'h29A7] = 8'h00;
RAM[16'h29A8] = 8'h00;
RAM[16'h29A9] = 8'h00;
RAM[16'h29AA] = 8'h00;
RAM[16'h29AB] = 8'h00;
RAM[16'h29AC] = 8'h00;
RAM[16'h29AD] = 8'h00;
RAM[16'h29AE] = 8'h00;
RAM[16'h29AF] = 8'h00;
RAM[16'h29B0] = 8'h00;
RAM[16'h29B1] = 8'h00;
RAM[16'h29B2] = 8'h00;
RAM[16'h29B3] = 8'h00;
RAM[16'h29B4] = 8'h00;
RAM[16'h29B5] = 8'h00;
RAM[16'h29B6] = 8'h00;
RAM[16'h29B7] = 8'h00;
RAM[16'h29B8] = 8'h00;
RAM[16'h29B9] = 8'h00;
RAM[16'h29BA] = 8'h00;
RAM[16'h29BB] = 8'h00;
RAM[16'h29BC] = 8'h00;
RAM[16'h29BD] = 8'h00;
RAM[16'h29BE] = 8'h00;
RAM[16'h29BF] = 8'h00;
RAM[16'h29C0] = 8'h00;
RAM[16'h29C1] = 8'h00;
RAM[16'h29C2] = 8'h00;
RAM[16'h29C3] = 8'h00;
RAM[16'h29C4] = 8'h00;
RAM[16'h29C5] = 8'h00;
RAM[16'h29C6] = 8'h00;
RAM[16'h29C7] = 8'h00;
RAM[16'h29C8] = 8'h00;
RAM[16'h29C9] = 8'h00;
RAM[16'h29CA] = 8'h00;
RAM[16'h29CB] = 8'h00;
RAM[16'h29CC] = 8'h00;
RAM[16'h29CD] = 8'h00;
RAM[16'h29CE] = 8'h00;
RAM[16'h29CF] = 8'h00;
RAM[16'h29D0] = 8'h00;
RAM[16'h29D1] = 8'h00;
RAM[16'h29D2] = 8'h00;
RAM[16'h29D3] = 8'h00;
RAM[16'h29D4] = 8'h00;
RAM[16'h29D5] = 8'h00;
RAM[16'h29D6] = 8'h00;
RAM[16'h29D7] = 8'h00;
RAM[16'h29D8] = 8'h00;
RAM[16'h29D9] = 8'h00;
RAM[16'h29DA] = 8'h00;
RAM[16'h29DB] = 8'h00;
RAM[16'h29DC] = 8'h00;
RAM[16'h29DD] = 8'h00;
RAM[16'h29DE] = 8'h00;
RAM[16'h29DF] = 8'h00;
RAM[16'h29E0] = 8'h00;
RAM[16'h29E1] = 8'h00;
RAM[16'h29E2] = 8'h00;
RAM[16'h29E3] = 8'h00;
RAM[16'h29E4] = 8'h00;
RAM[16'h29E5] = 8'h00;
RAM[16'h29E6] = 8'h00;
RAM[16'h29E7] = 8'h00;
RAM[16'h29E8] = 8'h00;
RAM[16'h29E9] = 8'h00;
RAM[16'h29EA] = 8'h00;
RAM[16'h29EB] = 8'h00;
RAM[16'h29EC] = 8'h00;
RAM[16'h29ED] = 8'h00;
RAM[16'h29EE] = 8'h00;
RAM[16'h29EF] = 8'h00;
RAM[16'h29F0] = 8'h00;
RAM[16'h29F1] = 8'h00;
RAM[16'h29F2] = 8'h00;
RAM[16'h29F3] = 8'h00;
RAM[16'h29F4] = 8'h00;
RAM[16'h29F5] = 8'h00;
RAM[16'h29F6] = 8'h00;
RAM[16'h29F7] = 8'h00;
RAM[16'h29F8] = 8'h00;
RAM[16'h29F9] = 8'h00;
RAM[16'h29FA] = 8'h00;
RAM[16'h29FB] = 8'h00;
RAM[16'h29FC] = 8'h00;
RAM[16'h29FD] = 8'h00;
RAM[16'h29FE] = 8'h00;
RAM[16'h29FF] = 8'h00;
RAM[16'h2A00] = 8'h00;
RAM[16'h2A01] = 8'h00;
RAM[16'h2A02] = 8'h00;
RAM[16'h2A03] = 8'h00;
RAM[16'h2A04] = 8'h00;
RAM[16'h2A05] = 8'h00;
RAM[16'h2A06] = 8'h00;
RAM[16'h2A07] = 8'h00;
RAM[16'h2A08] = 8'h00;
RAM[16'h2A09] = 8'h00;
RAM[16'h2A0A] = 8'h00;
RAM[16'h2A0B] = 8'h00;
RAM[16'h2A0C] = 8'h00;
RAM[16'h2A0D] = 8'h00;
RAM[16'h2A0E] = 8'h00;
RAM[16'h2A0F] = 8'h00;
RAM[16'h2A10] = 8'h00;
RAM[16'h2A11] = 8'h00;
RAM[16'h2A12] = 8'h00;
RAM[16'h2A13] = 8'h00;
RAM[16'h2A14] = 8'h00;
RAM[16'h2A15] = 8'h00;
RAM[16'h2A16] = 8'h00;
RAM[16'h2A17] = 8'h00;
RAM[16'h2A18] = 8'h00;
RAM[16'h2A19] = 8'h00;
RAM[16'h2A1A] = 8'h00;
RAM[16'h2A1B] = 8'h00;
RAM[16'h2A1C] = 8'h00;
RAM[16'h2A1D] = 8'h00;
RAM[16'h2A1E] = 8'h00;
RAM[16'h2A1F] = 8'h00;
RAM[16'h2A20] = 8'h00;
RAM[16'h2A21] = 8'h00;
RAM[16'h2A22] = 8'h00;
RAM[16'h2A23] = 8'h00;
RAM[16'h2A24] = 8'h00;
RAM[16'h2A25] = 8'h00;
RAM[16'h2A26] = 8'h00;
RAM[16'h2A27] = 8'h00;
RAM[16'h2A28] = 8'h00;
RAM[16'h2A29] = 8'h00;
RAM[16'h2A2A] = 8'h00;
RAM[16'h2A2B] = 8'h00;
RAM[16'h2A2C] = 8'h00;
RAM[16'h2A2D] = 8'h00;
RAM[16'h2A2E] = 8'h00;
RAM[16'h2A2F] = 8'h00;
RAM[16'h2A30] = 8'h00;
RAM[16'h2A31] = 8'h00;
RAM[16'h2A32] = 8'h00;
RAM[16'h2A33] = 8'h00;
RAM[16'h2A34] = 8'h00;
RAM[16'h2A35] = 8'h00;
RAM[16'h2A36] = 8'h00;
RAM[16'h2A37] = 8'h00;
RAM[16'h2A38] = 8'h00;
RAM[16'h2A39] = 8'h00;
RAM[16'h2A3A] = 8'h00;
RAM[16'h2A3B] = 8'h00;
RAM[16'h2A3C] = 8'h00;
RAM[16'h2A3D] = 8'h00;
RAM[16'h2A3E] = 8'h00;
RAM[16'h2A3F] = 8'h00;
RAM[16'h2A40] = 8'h00;
RAM[16'h2A41] = 8'h00;
RAM[16'h2A42] = 8'h00;
RAM[16'h2A43] = 8'h00;
RAM[16'h2A44] = 8'h00;
RAM[16'h2A45] = 8'h00;
RAM[16'h2A46] = 8'h00;
RAM[16'h2A47] = 8'h00;
RAM[16'h2A48] = 8'h00;
RAM[16'h2A49] = 8'h00;
RAM[16'h2A4A] = 8'h00;
RAM[16'h2A4B] = 8'h00;
RAM[16'h2A4C] = 8'h00;
RAM[16'h2A4D] = 8'h00;
RAM[16'h2A4E] = 8'h00;
RAM[16'h2A4F] = 8'h00;
RAM[16'h2A50] = 8'h00;
RAM[16'h2A51] = 8'h00;
RAM[16'h2A52] = 8'h00;
RAM[16'h2A53] = 8'h00;
RAM[16'h2A54] = 8'h00;
RAM[16'h2A55] = 8'h00;
RAM[16'h2A56] = 8'h00;
RAM[16'h2A57] = 8'h00;
RAM[16'h2A58] = 8'h00;
RAM[16'h2A59] = 8'h00;
RAM[16'h2A5A] = 8'h00;
RAM[16'h2A5B] = 8'h00;
RAM[16'h2A5C] = 8'h00;
RAM[16'h2A5D] = 8'h00;
RAM[16'h2A5E] = 8'h00;
RAM[16'h2A5F] = 8'h00;
RAM[16'h2A60] = 8'h00;
RAM[16'h2A61] = 8'h00;
RAM[16'h2A62] = 8'h00;
RAM[16'h2A63] = 8'h00;
RAM[16'h2A64] = 8'h00;
RAM[16'h2A65] = 8'h00;
RAM[16'h2A66] = 8'h00;
RAM[16'h2A67] = 8'h00;
RAM[16'h2A68] = 8'h00;
RAM[16'h2A69] = 8'h00;
RAM[16'h2A6A] = 8'h00;
RAM[16'h2A6B] = 8'h00;
RAM[16'h2A6C] = 8'h00;
RAM[16'h2A6D] = 8'h00;
RAM[16'h2A6E] = 8'h00;
RAM[16'h2A6F] = 8'h00;
RAM[16'h2A70] = 8'h00;
RAM[16'h2A71] = 8'h00;
RAM[16'h2A72] = 8'h00;
RAM[16'h2A73] = 8'h00;
RAM[16'h2A74] = 8'h00;
RAM[16'h2A75] = 8'h00;
RAM[16'h2A76] = 8'h00;
RAM[16'h2A77] = 8'h00;
RAM[16'h2A78] = 8'h00;
RAM[16'h2A79] = 8'h00;
RAM[16'h2A7A] = 8'h00;
RAM[16'h2A7B] = 8'h00;
RAM[16'h2A7C] = 8'h00;
RAM[16'h2A7D] = 8'h00;
RAM[16'h2A7E] = 8'h00;
RAM[16'h2A7F] = 8'h00;
RAM[16'h2A80] = 8'h00;
RAM[16'h2A81] = 8'h00;
RAM[16'h2A82] = 8'h00;
RAM[16'h2A83] = 8'h00;
RAM[16'h2A84] = 8'h00;
RAM[16'h2A85] = 8'h00;
RAM[16'h2A86] = 8'h00;
RAM[16'h2A87] = 8'h00;
RAM[16'h2A88] = 8'h00;
RAM[16'h2A89] = 8'h00;
RAM[16'h2A8A] = 8'h00;
RAM[16'h2A8B] = 8'h00;
RAM[16'h2A8C] = 8'h00;
RAM[16'h2A8D] = 8'h00;
RAM[16'h2A8E] = 8'h00;
RAM[16'h2A8F] = 8'h00;
RAM[16'h2A90] = 8'h00;
RAM[16'h2A91] = 8'h00;
RAM[16'h2A92] = 8'h00;
RAM[16'h2A93] = 8'h00;
RAM[16'h2A94] = 8'h00;
RAM[16'h2A95] = 8'h00;
RAM[16'h2A96] = 8'h00;
RAM[16'h2A97] = 8'h00;
RAM[16'h2A98] = 8'h00;
RAM[16'h2A99] = 8'h00;
RAM[16'h2A9A] = 8'h00;
RAM[16'h2A9B] = 8'h00;
RAM[16'h2A9C] = 8'h00;
RAM[16'h2A9D] = 8'h00;
RAM[16'h2A9E] = 8'h00;
RAM[16'h2A9F] = 8'h00;
RAM[16'h2AA0] = 8'h00;
RAM[16'h2AA1] = 8'h00;
RAM[16'h2AA2] = 8'h00;
RAM[16'h2AA3] = 8'h00;
RAM[16'h2AA4] = 8'h00;
RAM[16'h2AA5] = 8'h00;
RAM[16'h2AA6] = 8'h00;
RAM[16'h2AA7] = 8'h00;
RAM[16'h2AA8] = 8'h00;
RAM[16'h2AA9] = 8'h00;
RAM[16'h2AAA] = 8'h00;
RAM[16'h2AAB] = 8'h00;
RAM[16'h2AAC] = 8'h00;
RAM[16'h2AAD] = 8'h00;
RAM[16'h2AAE] = 8'h00;
RAM[16'h2AAF] = 8'h00;
RAM[16'h2AB0] = 8'h00;
RAM[16'h2AB1] = 8'h00;
RAM[16'h2AB2] = 8'h00;
RAM[16'h2AB3] = 8'h00;
RAM[16'h2AB4] = 8'h00;
RAM[16'h2AB5] = 8'h00;
RAM[16'h2AB6] = 8'h00;
RAM[16'h2AB7] = 8'h00;
RAM[16'h2AB8] = 8'h00;
RAM[16'h2AB9] = 8'h00;
RAM[16'h2ABA] = 8'h00;
RAM[16'h2ABB] = 8'h00;
RAM[16'h2ABC] = 8'h00;
RAM[16'h2ABD] = 8'h00;
RAM[16'h2ABE] = 8'h00;
RAM[16'h2ABF] = 8'h00;
RAM[16'h2AC0] = 8'h00;
RAM[16'h2AC1] = 8'h00;
RAM[16'h2AC2] = 8'h00;
RAM[16'h2AC3] = 8'h00;
RAM[16'h2AC4] = 8'h00;
RAM[16'h2AC5] = 8'h00;
RAM[16'h2AC6] = 8'h00;
RAM[16'h2AC7] = 8'h00;
RAM[16'h2AC8] = 8'h00;
RAM[16'h2AC9] = 8'h00;
RAM[16'h2ACA] = 8'h00;
RAM[16'h2ACB] = 8'h00;
RAM[16'h2ACC] = 8'h00;
RAM[16'h2ACD] = 8'h00;
RAM[16'h2ACE] = 8'h00;
RAM[16'h2ACF] = 8'h00;
RAM[16'h2AD0] = 8'h00;
RAM[16'h2AD1] = 8'h00;
RAM[16'h2AD2] = 8'h00;
RAM[16'h2AD3] = 8'h00;
RAM[16'h2AD4] = 8'h00;
RAM[16'h2AD5] = 8'h00;
RAM[16'h2AD6] = 8'h00;
RAM[16'h2AD7] = 8'h00;
RAM[16'h2AD8] = 8'h00;
RAM[16'h2AD9] = 8'h00;
RAM[16'h2ADA] = 8'h00;
RAM[16'h2ADB] = 8'h00;
RAM[16'h2ADC] = 8'h00;
RAM[16'h2ADD] = 8'h00;
RAM[16'h2ADE] = 8'h00;
RAM[16'h2ADF] = 8'h00;
RAM[16'h2AE0] = 8'h00;
RAM[16'h2AE1] = 8'h00;
RAM[16'h2AE2] = 8'h00;
RAM[16'h2AE3] = 8'h00;
RAM[16'h2AE4] = 8'h00;
RAM[16'h2AE5] = 8'h00;
RAM[16'h2AE6] = 8'h00;
RAM[16'h2AE7] = 8'h00;
RAM[16'h2AE8] = 8'h00;
RAM[16'h2AE9] = 8'h00;
RAM[16'h2AEA] = 8'h00;
RAM[16'h2AEB] = 8'h00;
RAM[16'h2AEC] = 8'h00;
RAM[16'h2AED] = 8'h00;
RAM[16'h2AEE] = 8'h00;
RAM[16'h2AEF] = 8'h00;
RAM[16'h2AF0] = 8'h00;
RAM[16'h2AF1] = 8'h00;
RAM[16'h2AF2] = 8'h00;
RAM[16'h2AF3] = 8'h00;
RAM[16'h2AF4] = 8'h00;
RAM[16'h2AF5] = 8'h00;
RAM[16'h2AF6] = 8'h00;
RAM[16'h2AF7] = 8'h00;
RAM[16'h2AF8] = 8'h00;
RAM[16'h2AF9] = 8'h00;
RAM[16'h2AFA] = 8'h00;
RAM[16'h2AFB] = 8'h00;
RAM[16'h2AFC] = 8'h00;
RAM[16'h2AFD] = 8'h00;
RAM[16'h2AFE] = 8'h00;
RAM[16'h2AFF] = 8'h00;
RAM[16'h2B00] = 8'h00;
RAM[16'h2B01] = 8'h00;
RAM[16'h2B02] = 8'h00;
RAM[16'h2B03] = 8'h00;
RAM[16'h2B04] = 8'h00;
RAM[16'h2B05] = 8'h00;
RAM[16'h2B06] = 8'h00;
RAM[16'h2B07] = 8'h00;
RAM[16'h2B08] = 8'h00;
RAM[16'h2B09] = 8'h00;
RAM[16'h2B0A] = 8'h00;
RAM[16'h2B0B] = 8'h00;
RAM[16'h2B0C] = 8'h00;
RAM[16'h2B0D] = 8'h00;
RAM[16'h2B0E] = 8'h00;
RAM[16'h2B0F] = 8'h00;
RAM[16'h2B10] = 8'h00;
RAM[16'h2B11] = 8'h00;
RAM[16'h2B12] = 8'h00;
RAM[16'h2B13] = 8'h00;
RAM[16'h2B14] = 8'h00;
RAM[16'h2B15] = 8'h00;
RAM[16'h2B16] = 8'h00;
RAM[16'h2B17] = 8'h00;
RAM[16'h2B18] = 8'h00;
RAM[16'h2B19] = 8'h00;
RAM[16'h2B1A] = 8'h00;
RAM[16'h2B1B] = 8'h00;
RAM[16'h2B1C] = 8'h00;
RAM[16'h2B1D] = 8'h00;
RAM[16'h2B1E] = 8'h00;
RAM[16'h2B1F] = 8'h00;
RAM[16'h2B20] = 8'h00;
RAM[16'h2B21] = 8'h00;
RAM[16'h2B22] = 8'h00;
RAM[16'h2B23] = 8'h00;
RAM[16'h2B24] = 8'h00;
RAM[16'h2B25] = 8'h00;
RAM[16'h2B26] = 8'h00;
RAM[16'h2B27] = 8'h00;
RAM[16'h2B28] = 8'h00;
RAM[16'h2B29] = 8'h00;
RAM[16'h2B2A] = 8'h00;
RAM[16'h2B2B] = 8'h00;
RAM[16'h2B2C] = 8'h00;
RAM[16'h2B2D] = 8'h00;
RAM[16'h2B2E] = 8'h00;
RAM[16'h2B2F] = 8'h00;
RAM[16'h2B30] = 8'h00;
RAM[16'h2B31] = 8'h00;
RAM[16'h2B32] = 8'h00;
RAM[16'h2B33] = 8'h00;
RAM[16'h2B34] = 8'h00;
RAM[16'h2B35] = 8'h00;
RAM[16'h2B36] = 8'h00;
RAM[16'h2B37] = 8'h00;
RAM[16'h2B38] = 8'h00;
RAM[16'h2B39] = 8'h00;
RAM[16'h2B3A] = 8'h00;
RAM[16'h2B3B] = 8'h00;
RAM[16'h2B3C] = 8'h00;
RAM[16'h2B3D] = 8'h00;
RAM[16'h2B3E] = 8'h00;
RAM[16'h2B3F] = 8'h00;
RAM[16'h2B40] = 8'h00;
RAM[16'h2B41] = 8'h00;
RAM[16'h2B42] = 8'h00;
RAM[16'h2B43] = 8'h00;
RAM[16'h2B44] = 8'h00;
RAM[16'h2B45] = 8'h00;
RAM[16'h2B46] = 8'h00;
RAM[16'h2B47] = 8'h00;
RAM[16'h2B48] = 8'h00;
RAM[16'h2B49] = 8'h00;
RAM[16'h2B4A] = 8'h00;
RAM[16'h2B4B] = 8'h00;
RAM[16'h2B4C] = 8'h00;
RAM[16'h2B4D] = 8'h00;
RAM[16'h2B4E] = 8'h00;
RAM[16'h2B4F] = 8'h00;
RAM[16'h2B50] = 8'h00;
RAM[16'h2B51] = 8'h00;
RAM[16'h2B52] = 8'h00;
RAM[16'h2B53] = 8'h00;
RAM[16'h2B54] = 8'h00;
RAM[16'h2B55] = 8'h00;
RAM[16'h2B56] = 8'h00;
RAM[16'h2B57] = 8'h00;
RAM[16'h2B58] = 8'h00;
RAM[16'h2B59] = 8'h00;
RAM[16'h2B5A] = 8'h00;
RAM[16'h2B5B] = 8'h00;
RAM[16'h2B5C] = 8'h00;
RAM[16'h2B5D] = 8'h00;
RAM[16'h2B5E] = 8'h00;
RAM[16'h2B5F] = 8'h00;
RAM[16'h2B60] = 8'h00;
RAM[16'h2B61] = 8'h00;
RAM[16'h2B62] = 8'h00;
RAM[16'h2B63] = 8'h00;
RAM[16'h2B64] = 8'h00;
RAM[16'h2B65] = 8'h00;
RAM[16'h2B66] = 8'h00;
RAM[16'h2B67] = 8'h00;
RAM[16'h2B68] = 8'h00;
RAM[16'h2B69] = 8'h00;
RAM[16'h2B6A] = 8'h00;
RAM[16'h2B6B] = 8'h00;
RAM[16'h2B6C] = 8'h00;
RAM[16'h2B6D] = 8'h00;
RAM[16'h2B6E] = 8'h00;
RAM[16'h2B6F] = 8'h00;
RAM[16'h2B70] = 8'h00;
RAM[16'h2B71] = 8'h00;
RAM[16'h2B72] = 8'h00;
RAM[16'h2B73] = 8'h00;
RAM[16'h2B74] = 8'h00;
RAM[16'h2B75] = 8'h00;
RAM[16'h2B76] = 8'h00;
RAM[16'h2B77] = 8'h00;
RAM[16'h2B78] = 8'h00;
RAM[16'h2B79] = 8'h00;
RAM[16'h2B7A] = 8'h00;
RAM[16'h2B7B] = 8'h00;
RAM[16'h2B7C] = 8'h00;
RAM[16'h2B7D] = 8'h00;
RAM[16'h2B7E] = 8'h00;
RAM[16'h2B7F] = 8'h00;
RAM[16'h2B80] = 8'h00;
RAM[16'h2B81] = 8'h00;
RAM[16'h2B82] = 8'h00;
RAM[16'h2B83] = 8'h00;
RAM[16'h2B84] = 8'h00;
RAM[16'h2B85] = 8'h00;
RAM[16'h2B86] = 8'h00;
RAM[16'h2B87] = 8'h00;
RAM[16'h2B88] = 8'h00;
RAM[16'h2B89] = 8'h00;
RAM[16'h2B8A] = 8'h00;
RAM[16'h2B8B] = 8'h00;
RAM[16'h2B8C] = 8'h00;
RAM[16'h2B8D] = 8'h00;
RAM[16'h2B8E] = 8'h00;
RAM[16'h2B8F] = 8'h00;
RAM[16'h2B90] = 8'h00;
RAM[16'h2B91] = 8'h00;
RAM[16'h2B92] = 8'h00;
RAM[16'h2B93] = 8'h00;
RAM[16'h2B94] = 8'h00;
RAM[16'h2B95] = 8'h00;
RAM[16'h2B96] = 8'h00;
RAM[16'h2B97] = 8'h00;
RAM[16'h2B98] = 8'h00;
RAM[16'h2B99] = 8'h00;
RAM[16'h2B9A] = 8'h00;
RAM[16'h2B9B] = 8'h00;
RAM[16'h2B9C] = 8'h00;
RAM[16'h2B9D] = 8'h00;
RAM[16'h2B9E] = 8'h00;
RAM[16'h2B9F] = 8'h00;
RAM[16'h2BA0] = 8'h00;
RAM[16'h2BA1] = 8'h00;
RAM[16'h2BA2] = 8'h00;
RAM[16'h2BA3] = 8'h00;
RAM[16'h2BA4] = 8'h00;
RAM[16'h2BA5] = 8'h00;
RAM[16'h2BA6] = 8'h00;
RAM[16'h2BA7] = 8'h00;
RAM[16'h2BA8] = 8'h00;
RAM[16'h2BA9] = 8'h00;
RAM[16'h2BAA] = 8'h00;
RAM[16'h2BAB] = 8'h00;
RAM[16'h2BAC] = 8'h00;
RAM[16'h2BAD] = 8'h00;
RAM[16'h2BAE] = 8'h00;
RAM[16'h2BAF] = 8'h00;
RAM[16'h2BB0] = 8'h00;
RAM[16'h2BB1] = 8'h00;
RAM[16'h2BB2] = 8'h00;
RAM[16'h2BB3] = 8'h00;
RAM[16'h2BB4] = 8'h00;
RAM[16'h2BB5] = 8'h00;
RAM[16'h2BB6] = 8'h00;
RAM[16'h2BB7] = 8'h00;
RAM[16'h2BB8] = 8'h00;
RAM[16'h2BB9] = 8'h00;
RAM[16'h2BBA] = 8'h00;
RAM[16'h2BBB] = 8'h00;
RAM[16'h2BBC] = 8'h00;
RAM[16'h2BBD] = 8'h00;
RAM[16'h2BBE] = 8'h00;
RAM[16'h2BBF] = 8'h00;
RAM[16'h2BC0] = 8'h00;
RAM[16'h2BC1] = 8'h00;
RAM[16'h2BC2] = 8'h00;
RAM[16'h2BC3] = 8'h00;
RAM[16'h2BC4] = 8'h00;
RAM[16'h2BC5] = 8'h00;
RAM[16'h2BC6] = 8'h00;
RAM[16'h2BC7] = 8'h00;
RAM[16'h2BC8] = 8'h00;
RAM[16'h2BC9] = 8'h00;
RAM[16'h2BCA] = 8'h00;
RAM[16'h2BCB] = 8'h00;
RAM[16'h2BCC] = 8'h00;
RAM[16'h2BCD] = 8'h00;
RAM[16'h2BCE] = 8'h00;
RAM[16'h2BCF] = 8'h00;
RAM[16'h2BD0] = 8'h00;
RAM[16'h2BD1] = 8'h00;
RAM[16'h2BD2] = 8'h00;
RAM[16'h2BD3] = 8'h00;
RAM[16'h2BD4] = 8'h00;
RAM[16'h2BD5] = 8'h00;
RAM[16'h2BD6] = 8'h00;
RAM[16'h2BD7] = 8'h00;
RAM[16'h2BD8] = 8'h00;
RAM[16'h2BD9] = 8'h00;
RAM[16'h2BDA] = 8'h00;
RAM[16'h2BDB] = 8'h00;
RAM[16'h2BDC] = 8'h00;
RAM[16'h2BDD] = 8'h00;
RAM[16'h2BDE] = 8'h00;
RAM[16'h2BDF] = 8'h00;
RAM[16'h2BE0] = 8'h00;
RAM[16'h2BE1] = 8'h00;
RAM[16'h2BE2] = 8'h00;
RAM[16'h2BE3] = 8'h00;
RAM[16'h2BE4] = 8'h00;
RAM[16'h2BE5] = 8'h00;
RAM[16'h2BE6] = 8'h00;
RAM[16'h2BE7] = 8'h00;
RAM[16'h2BE8] = 8'h00;
RAM[16'h2BE9] = 8'h00;
RAM[16'h2BEA] = 8'h00;
RAM[16'h2BEB] = 8'h00;
RAM[16'h2BEC] = 8'h00;
RAM[16'h2BED] = 8'h00;
RAM[16'h2BEE] = 8'h00;
RAM[16'h2BEF] = 8'h00;
RAM[16'h2BF0] = 8'h00;
RAM[16'h2BF1] = 8'h00;
RAM[16'h2BF2] = 8'h00;
RAM[16'h2BF3] = 8'h00;
RAM[16'h2BF4] = 8'h00;
RAM[16'h2BF5] = 8'h00;
RAM[16'h2BF6] = 8'h00;
RAM[16'h2BF7] = 8'h00;
RAM[16'h2BF8] = 8'h00;
RAM[16'h2BF9] = 8'h00;
RAM[16'h2BFA] = 8'h00;
RAM[16'h2BFB] = 8'h00;
RAM[16'h2BFC] = 8'h00;
RAM[16'h2BFD] = 8'h00;
RAM[16'h2BFE] = 8'h00;
RAM[16'h2BFF] = 8'h00;
RAM[16'h2C00] = 8'h00;
RAM[16'h2C01] = 8'h00;
RAM[16'h2C02] = 8'h00;
RAM[16'h2C03] = 8'h00;
RAM[16'h2C04] = 8'h00;
RAM[16'h2C05] = 8'h00;
RAM[16'h2C06] = 8'h00;
RAM[16'h2C07] = 8'h00;
RAM[16'h2C08] = 8'h00;
RAM[16'h2C09] = 8'h00;
RAM[16'h2C0A] = 8'h00;
RAM[16'h2C0B] = 8'h00;
RAM[16'h2C0C] = 8'h00;
RAM[16'h2C0D] = 8'h00;
RAM[16'h2C0E] = 8'h00;
RAM[16'h2C0F] = 8'h00;
RAM[16'h2C10] = 8'h00;
RAM[16'h2C11] = 8'h00;
RAM[16'h2C12] = 8'h00;
RAM[16'h2C13] = 8'h00;
RAM[16'h2C14] = 8'h00;
RAM[16'h2C15] = 8'h00;
RAM[16'h2C16] = 8'h00;
RAM[16'h2C17] = 8'h00;
RAM[16'h2C18] = 8'h00;
RAM[16'h2C19] = 8'h00;
RAM[16'h2C1A] = 8'h00;
RAM[16'h2C1B] = 8'h00;
RAM[16'h2C1C] = 8'h00;
RAM[16'h2C1D] = 8'h00;
RAM[16'h2C1E] = 8'h00;
RAM[16'h2C1F] = 8'h00;
RAM[16'h2C20] = 8'h00;
RAM[16'h2C21] = 8'h00;
RAM[16'h2C22] = 8'h00;
RAM[16'h2C23] = 8'h00;
RAM[16'h2C24] = 8'h00;
RAM[16'h2C25] = 8'h00;
RAM[16'h2C26] = 8'h00;
RAM[16'h2C27] = 8'h00;
RAM[16'h2C28] = 8'h00;
RAM[16'h2C29] = 8'h00;
RAM[16'h2C2A] = 8'h00;
RAM[16'h2C2B] = 8'h00;
RAM[16'h2C2C] = 8'h00;
RAM[16'h2C2D] = 8'h00;
RAM[16'h2C2E] = 8'h00;
RAM[16'h2C2F] = 8'h00;
RAM[16'h2C30] = 8'h00;
RAM[16'h2C31] = 8'h00;
RAM[16'h2C32] = 8'h00;
RAM[16'h2C33] = 8'h00;
RAM[16'h2C34] = 8'h00;
RAM[16'h2C35] = 8'h00;
RAM[16'h2C36] = 8'h00;
RAM[16'h2C37] = 8'h00;
RAM[16'h2C38] = 8'h00;
RAM[16'h2C39] = 8'h00;
RAM[16'h2C3A] = 8'h00;
RAM[16'h2C3B] = 8'h00;
RAM[16'h2C3C] = 8'h00;
RAM[16'h2C3D] = 8'h00;
RAM[16'h2C3E] = 8'h00;
RAM[16'h2C3F] = 8'h00;
RAM[16'h2C40] = 8'h00;
RAM[16'h2C41] = 8'h00;
RAM[16'h2C42] = 8'h00;
RAM[16'h2C43] = 8'h00;
RAM[16'h2C44] = 8'h00;
RAM[16'h2C45] = 8'h00;
RAM[16'h2C46] = 8'h00;
RAM[16'h2C47] = 8'h00;
RAM[16'h2C48] = 8'h00;
RAM[16'h2C49] = 8'h00;
RAM[16'h2C4A] = 8'h00;
RAM[16'h2C4B] = 8'h00;
RAM[16'h2C4C] = 8'h00;
RAM[16'h2C4D] = 8'h00;
RAM[16'h2C4E] = 8'h00;
RAM[16'h2C4F] = 8'h00;
RAM[16'h2C50] = 8'h00;
RAM[16'h2C51] = 8'h00;
RAM[16'h2C52] = 8'h00;
RAM[16'h2C53] = 8'h00;
RAM[16'h2C54] = 8'h00;
RAM[16'h2C55] = 8'h00;
RAM[16'h2C56] = 8'h00;
RAM[16'h2C57] = 8'h00;
RAM[16'h2C58] = 8'h00;
RAM[16'h2C59] = 8'h00;
RAM[16'h2C5A] = 8'h00;
RAM[16'h2C5B] = 8'h00;
RAM[16'h2C5C] = 8'h00;
RAM[16'h2C5D] = 8'h00;
RAM[16'h2C5E] = 8'h00;
RAM[16'h2C5F] = 8'h00;
RAM[16'h2C60] = 8'h00;
RAM[16'h2C61] = 8'h00;
RAM[16'h2C62] = 8'h00;
RAM[16'h2C63] = 8'h00;
RAM[16'h2C64] = 8'h00;
RAM[16'h2C65] = 8'h00;
RAM[16'h2C66] = 8'h00;
RAM[16'h2C67] = 8'h00;
RAM[16'h2C68] = 8'h00;
RAM[16'h2C69] = 8'h00;
RAM[16'h2C6A] = 8'h00;
RAM[16'h2C6B] = 8'h00;
RAM[16'h2C6C] = 8'h00;
RAM[16'h2C6D] = 8'h00;
RAM[16'h2C6E] = 8'h00;
RAM[16'h2C6F] = 8'h00;
RAM[16'h2C70] = 8'h00;
RAM[16'h2C71] = 8'h00;
RAM[16'h2C72] = 8'h00;
RAM[16'h2C73] = 8'h00;
RAM[16'h2C74] = 8'h00;
RAM[16'h2C75] = 8'h00;
RAM[16'h2C76] = 8'h00;
RAM[16'h2C77] = 8'h00;
RAM[16'h2C78] = 8'h00;
RAM[16'h2C79] = 8'h00;
RAM[16'h2C7A] = 8'h00;
RAM[16'h2C7B] = 8'h00;
RAM[16'h2C7C] = 8'h00;
RAM[16'h2C7D] = 8'h00;
RAM[16'h2C7E] = 8'h00;
RAM[16'h2C7F] = 8'h00;
RAM[16'h2C80] = 8'h00;
RAM[16'h2C81] = 8'h00;
RAM[16'h2C82] = 8'h00;
RAM[16'h2C83] = 8'h00;
RAM[16'h2C84] = 8'h00;
RAM[16'h2C85] = 8'h00;
RAM[16'h2C86] = 8'h00;
RAM[16'h2C87] = 8'h00;
RAM[16'h2C88] = 8'h00;
RAM[16'h2C89] = 8'h00;
RAM[16'h2C8A] = 8'h00;
RAM[16'h2C8B] = 8'h00;
RAM[16'h2C8C] = 8'h00;
RAM[16'h2C8D] = 8'h00;
RAM[16'h2C8E] = 8'h00;
RAM[16'h2C8F] = 8'h00;
RAM[16'h2C90] = 8'h00;
RAM[16'h2C91] = 8'h00;
RAM[16'h2C92] = 8'h00;
RAM[16'h2C93] = 8'h00;
RAM[16'h2C94] = 8'h00;
RAM[16'h2C95] = 8'h00;
RAM[16'h2C96] = 8'h00;
RAM[16'h2C97] = 8'h00;
RAM[16'h2C98] = 8'h00;
RAM[16'h2C99] = 8'h00;
RAM[16'h2C9A] = 8'h00;
RAM[16'h2C9B] = 8'h00;
RAM[16'h2C9C] = 8'h00;
RAM[16'h2C9D] = 8'h00;
RAM[16'h2C9E] = 8'h00;
RAM[16'h2C9F] = 8'h00;
RAM[16'h2CA0] = 8'h00;
RAM[16'h2CA1] = 8'h00;
RAM[16'h2CA2] = 8'h00;
RAM[16'h2CA3] = 8'h00;
RAM[16'h2CA4] = 8'h00;
RAM[16'h2CA5] = 8'h00;
RAM[16'h2CA6] = 8'h00;
RAM[16'h2CA7] = 8'h00;
RAM[16'h2CA8] = 8'h00;
RAM[16'h2CA9] = 8'h00;
RAM[16'h2CAA] = 8'h00;
RAM[16'h2CAB] = 8'h00;
RAM[16'h2CAC] = 8'h00;
RAM[16'h2CAD] = 8'h00;
RAM[16'h2CAE] = 8'h00;
RAM[16'h2CAF] = 8'h00;
RAM[16'h2CB0] = 8'h00;
RAM[16'h2CB1] = 8'h00;
RAM[16'h2CB2] = 8'h00;
RAM[16'h2CB3] = 8'h00;
RAM[16'h2CB4] = 8'h00;
RAM[16'h2CB5] = 8'h00;
RAM[16'h2CB6] = 8'h00;
RAM[16'h2CB7] = 8'h00;
RAM[16'h2CB8] = 8'h00;
RAM[16'h2CB9] = 8'h00;
RAM[16'h2CBA] = 8'h00;
RAM[16'h2CBB] = 8'h00;
RAM[16'h2CBC] = 8'h00;
RAM[16'h2CBD] = 8'h00;
RAM[16'h2CBE] = 8'h00;
RAM[16'h2CBF] = 8'h00;
RAM[16'h2CC0] = 8'h00;
RAM[16'h2CC1] = 8'h00;
RAM[16'h2CC2] = 8'h00;
RAM[16'h2CC3] = 8'h00;
RAM[16'h2CC4] = 8'h00;
RAM[16'h2CC5] = 8'h00;
RAM[16'h2CC6] = 8'h00;
RAM[16'h2CC7] = 8'h00;
RAM[16'h2CC8] = 8'h00;
RAM[16'h2CC9] = 8'h00;
RAM[16'h2CCA] = 8'h00;
RAM[16'h2CCB] = 8'h00;
RAM[16'h2CCC] = 8'h00;
RAM[16'h2CCD] = 8'h00;
RAM[16'h2CCE] = 8'h00;
RAM[16'h2CCF] = 8'h00;
RAM[16'h2CD0] = 8'h00;
RAM[16'h2CD1] = 8'h00;
RAM[16'h2CD2] = 8'h00;
RAM[16'h2CD3] = 8'h00;
RAM[16'h2CD4] = 8'h00;
RAM[16'h2CD5] = 8'h00;
RAM[16'h2CD6] = 8'h00;
RAM[16'h2CD7] = 8'h00;
RAM[16'h2CD8] = 8'h00;
RAM[16'h2CD9] = 8'h00;
RAM[16'h2CDA] = 8'h00;
RAM[16'h2CDB] = 8'h00;
RAM[16'h2CDC] = 8'h00;
RAM[16'h2CDD] = 8'h00;
RAM[16'h2CDE] = 8'h00;
RAM[16'h2CDF] = 8'h00;
RAM[16'h2CE0] = 8'h00;
RAM[16'h2CE1] = 8'h00;
RAM[16'h2CE2] = 8'h00;
RAM[16'h2CE3] = 8'h00;
RAM[16'h2CE4] = 8'h00;
RAM[16'h2CE5] = 8'h00;
RAM[16'h2CE6] = 8'h00;
RAM[16'h2CE7] = 8'h00;
RAM[16'h2CE8] = 8'h00;
RAM[16'h2CE9] = 8'h00;
RAM[16'h2CEA] = 8'h00;
RAM[16'h2CEB] = 8'h00;
RAM[16'h2CEC] = 8'h00;
RAM[16'h2CED] = 8'h00;
RAM[16'h2CEE] = 8'h00;
RAM[16'h2CEF] = 8'h00;
RAM[16'h2CF0] = 8'h00;
RAM[16'h2CF1] = 8'h00;
RAM[16'h2CF2] = 8'h00;
RAM[16'h2CF3] = 8'h00;
RAM[16'h2CF4] = 8'h00;
RAM[16'h2CF5] = 8'h00;
RAM[16'h2CF6] = 8'h00;
RAM[16'h2CF7] = 8'h00;
RAM[16'h2CF8] = 8'h00;
RAM[16'h2CF9] = 8'h00;
RAM[16'h2CFA] = 8'h00;
RAM[16'h2CFB] = 8'h00;
RAM[16'h2CFC] = 8'h00;
RAM[16'h2CFD] = 8'h00;
RAM[16'h2CFE] = 8'h00;
RAM[16'h2CFF] = 8'h00;
RAM[16'h2D00] = 8'h00;
RAM[16'h2D01] = 8'h00;
RAM[16'h2D02] = 8'h00;
RAM[16'h2D03] = 8'h00;
RAM[16'h2D04] = 8'h00;
RAM[16'h2D05] = 8'h00;
RAM[16'h2D06] = 8'h00;
RAM[16'h2D07] = 8'h00;
RAM[16'h2D08] = 8'h00;
RAM[16'h2D09] = 8'h00;
RAM[16'h2D0A] = 8'h00;
RAM[16'h2D0B] = 8'h00;
RAM[16'h2D0C] = 8'h00;
RAM[16'h2D0D] = 8'h00;
RAM[16'h2D0E] = 8'h00;
RAM[16'h2D0F] = 8'h00;
RAM[16'h2D10] = 8'h00;
RAM[16'h2D11] = 8'h00;
RAM[16'h2D12] = 8'h00;
RAM[16'h2D13] = 8'h00;
RAM[16'h2D14] = 8'h00;
RAM[16'h2D15] = 8'h00;
RAM[16'h2D16] = 8'h00;
RAM[16'h2D17] = 8'h00;
RAM[16'h2D18] = 8'h00;
RAM[16'h2D19] = 8'h00;
RAM[16'h2D1A] = 8'h00;
RAM[16'h2D1B] = 8'h00;
RAM[16'h2D1C] = 8'h00;
RAM[16'h2D1D] = 8'h00;
RAM[16'h2D1E] = 8'h00;
RAM[16'h2D1F] = 8'h00;
RAM[16'h2D20] = 8'h00;
RAM[16'h2D21] = 8'h00;
RAM[16'h2D22] = 8'h00;
RAM[16'h2D23] = 8'h00;
RAM[16'h2D24] = 8'h00;
RAM[16'h2D25] = 8'h00;
RAM[16'h2D26] = 8'h00;
RAM[16'h2D27] = 8'h00;
RAM[16'h2D28] = 8'h00;
RAM[16'h2D29] = 8'h00;
RAM[16'h2D2A] = 8'h00;
RAM[16'h2D2B] = 8'h00;
RAM[16'h2D2C] = 8'h00;
RAM[16'h2D2D] = 8'h00;
RAM[16'h2D2E] = 8'h00;
RAM[16'h2D2F] = 8'h00;
RAM[16'h2D30] = 8'h00;
RAM[16'h2D31] = 8'h00;
RAM[16'h2D32] = 8'h00;
RAM[16'h2D33] = 8'h00;
RAM[16'h2D34] = 8'h00;
RAM[16'h2D35] = 8'h00;
RAM[16'h2D36] = 8'h00;
RAM[16'h2D37] = 8'h00;
RAM[16'h2D38] = 8'h00;
RAM[16'h2D39] = 8'h00;
RAM[16'h2D3A] = 8'h00;
RAM[16'h2D3B] = 8'h00;
RAM[16'h2D3C] = 8'h00;
RAM[16'h2D3D] = 8'h00;
RAM[16'h2D3E] = 8'h00;
RAM[16'h2D3F] = 8'h00;
RAM[16'h2D40] = 8'h00;
RAM[16'h2D41] = 8'h00;
RAM[16'h2D42] = 8'h00;
RAM[16'h2D43] = 8'h00;
RAM[16'h2D44] = 8'h00;
RAM[16'h2D45] = 8'h00;
RAM[16'h2D46] = 8'h00;
RAM[16'h2D47] = 8'h00;
RAM[16'h2D48] = 8'h00;
RAM[16'h2D49] = 8'h00;
RAM[16'h2D4A] = 8'h00;
RAM[16'h2D4B] = 8'h00;
RAM[16'h2D4C] = 8'h00;
RAM[16'h2D4D] = 8'h00;
RAM[16'h2D4E] = 8'h00;
RAM[16'h2D4F] = 8'h00;
RAM[16'h2D50] = 8'h00;
RAM[16'h2D51] = 8'h00;
RAM[16'h2D52] = 8'h00;
RAM[16'h2D53] = 8'h00;
RAM[16'h2D54] = 8'h00;
RAM[16'h2D55] = 8'h00;
RAM[16'h2D56] = 8'h00;
RAM[16'h2D57] = 8'h00;
RAM[16'h2D58] = 8'h00;
RAM[16'h2D59] = 8'h00;
RAM[16'h2D5A] = 8'h00;
RAM[16'h2D5B] = 8'h00;
RAM[16'h2D5C] = 8'h00;
RAM[16'h2D5D] = 8'h00;
RAM[16'h2D5E] = 8'h00;
RAM[16'h2D5F] = 8'h00;
RAM[16'h2D60] = 8'h00;
RAM[16'h2D61] = 8'h00;
RAM[16'h2D62] = 8'h00;
RAM[16'h2D63] = 8'h00;
RAM[16'h2D64] = 8'h00;
RAM[16'h2D65] = 8'h00;
RAM[16'h2D66] = 8'h00;
RAM[16'h2D67] = 8'h00;
RAM[16'h2D68] = 8'h00;
RAM[16'h2D69] = 8'h00;
RAM[16'h2D6A] = 8'h00;
RAM[16'h2D6B] = 8'h00;
RAM[16'h2D6C] = 8'h00;
RAM[16'h2D6D] = 8'h00;
RAM[16'h2D6E] = 8'h00;
RAM[16'h2D6F] = 8'h00;
RAM[16'h2D70] = 8'h00;
RAM[16'h2D71] = 8'h00;
RAM[16'h2D72] = 8'h00;
RAM[16'h2D73] = 8'h00;
RAM[16'h2D74] = 8'h00;
RAM[16'h2D75] = 8'h00;
RAM[16'h2D76] = 8'h00;
RAM[16'h2D77] = 8'h00;
RAM[16'h2D78] = 8'h00;
RAM[16'h2D79] = 8'h00;
RAM[16'h2D7A] = 8'h00;
RAM[16'h2D7B] = 8'h00;
RAM[16'h2D7C] = 8'h00;
RAM[16'h2D7D] = 8'h00;
RAM[16'h2D7E] = 8'h00;
RAM[16'h2D7F] = 8'h00;
RAM[16'h2D80] = 8'h00;
RAM[16'h2D81] = 8'h00;
RAM[16'h2D82] = 8'h00;
RAM[16'h2D83] = 8'h00;
RAM[16'h2D84] = 8'h00;
RAM[16'h2D85] = 8'h00;
RAM[16'h2D86] = 8'h00;
RAM[16'h2D87] = 8'h00;
RAM[16'h2D88] = 8'h00;
RAM[16'h2D89] = 8'h00;
RAM[16'h2D8A] = 8'h00;
RAM[16'h2D8B] = 8'h00;
RAM[16'h2D8C] = 8'h00;
RAM[16'h2D8D] = 8'h00;
RAM[16'h2D8E] = 8'h00;
RAM[16'h2D8F] = 8'h00;
RAM[16'h2D90] = 8'h00;
RAM[16'h2D91] = 8'h00;
RAM[16'h2D92] = 8'h00;
RAM[16'h2D93] = 8'h00;
RAM[16'h2D94] = 8'h00;
RAM[16'h2D95] = 8'h00;
RAM[16'h2D96] = 8'h00;
RAM[16'h2D97] = 8'h00;
RAM[16'h2D98] = 8'h00;
RAM[16'h2D99] = 8'h00;
RAM[16'h2D9A] = 8'h00;
RAM[16'h2D9B] = 8'h00;
RAM[16'h2D9C] = 8'h00;
RAM[16'h2D9D] = 8'h00;
RAM[16'h2D9E] = 8'h00;
RAM[16'h2D9F] = 8'h00;
RAM[16'h2DA0] = 8'h00;
RAM[16'h2DA1] = 8'h00;
RAM[16'h2DA2] = 8'h00;
RAM[16'h2DA3] = 8'h00;
RAM[16'h2DA4] = 8'h00;
RAM[16'h2DA5] = 8'h00;
RAM[16'h2DA6] = 8'h00;
RAM[16'h2DA7] = 8'h00;
RAM[16'h2DA8] = 8'h00;
RAM[16'h2DA9] = 8'h00;
RAM[16'h2DAA] = 8'h00;
RAM[16'h2DAB] = 8'h00;
RAM[16'h2DAC] = 8'h00;
RAM[16'h2DAD] = 8'h00;
RAM[16'h2DAE] = 8'h00;
RAM[16'h2DAF] = 8'h00;
RAM[16'h2DB0] = 8'h00;
RAM[16'h2DB1] = 8'h00;
RAM[16'h2DB2] = 8'h00;
RAM[16'h2DB3] = 8'h00;
RAM[16'h2DB4] = 8'h00;
RAM[16'h2DB5] = 8'h00;
RAM[16'h2DB6] = 8'h00;
RAM[16'h2DB7] = 8'h00;
RAM[16'h2DB8] = 8'h00;
RAM[16'h2DB9] = 8'h00;
RAM[16'h2DBA] = 8'h00;
RAM[16'h2DBB] = 8'h00;
RAM[16'h2DBC] = 8'h00;
RAM[16'h2DBD] = 8'h00;
RAM[16'h2DBE] = 8'h00;
RAM[16'h2DBF] = 8'h00;
RAM[16'h2DC0] = 8'h00;
RAM[16'h2DC1] = 8'h00;
RAM[16'h2DC2] = 8'h00;
RAM[16'h2DC3] = 8'h00;
RAM[16'h2DC4] = 8'h00;
RAM[16'h2DC5] = 8'h00;
RAM[16'h2DC6] = 8'h00;
RAM[16'h2DC7] = 8'h00;
RAM[16'h2DC8] = 8'h00;
RAM[16'h2DC9] = 8'h00;
RAM[16'h2DCA] = 8'h00;
RAM[16'h2DCB] = 8'h00;
RAM[16'h2DCC] = 8'h00;
RAM[16'h2DCD] = 8'h00;
RAM[16'h2DCE] = 8'h00;
RAM[16'h2DCF] = 8'h00;
RAM[16'h2DD0] = 8'h00;
RAM[16'h2DD1] = 8'h00;
RAM[16'h2DD2] = 8'h00;
RAM[16'h2DD3] = 8'h00;
RAM[16'h2DD4] = 8'h00;
RAM[16'h2DD5] = 8'h00;
RAM[16'h2DD6] = 8'h00;
RAM[16'h2DD7] = 8'h00;
RAM[16'h2DD8] = 8'h00;
RAM[16'h2DD9] = 8'h00;
RAM[16'h2DDA] = 8'h00;
RAM[16'h2DDB] = 8'h00;
RAM[16'h2DDC] = 8'h00;
RAM[16'h2DDD] = 8'h00;
RAM[16'h2DDE] = 8'h00;
RAM[16'h2DDF] = 8'h00;
RAM[16'h2DE0] = 8'h00;
RAM[16'h2DE1] = 8'h00;
RAM[16'h2DE2] = 8'h00;
RAM[16'h2DE3] = 8'h00;
RAM[16'h2DE4] = 8'h00;
RAM[16'h2DE5] = 8'h00;
RAM[16'h2DE6] = 8'h00;
RAM[16'h2DE7] = 8'h00;
RAM[16'h2DE8] = 8'h00;
RAM[16'h2DE9] = 8'h00;
RAM[16'h2DEA] = 8'h00;
RAM[16'h2DEB] = 8'h00;
RAM[16'h2DEC] = 8'h00;
RAM[16'h2DED] = 8'h00;
RAM[16'h2DEE] = 8'h00;
RAM[16'h2DEF] = 8'h00;
RAM[16'h2DF0] = 8'h00;
RAM[16'h2DF1] = 8'h00;
RAM[16'h2DF2] = 8'h00;
RAM[16'h2DF3] = 8'h00;
RAM[16'h2DF4] = 8'h00;
RAM[16'h2DF5] = 8'h00;
RAM[16'h2DF6] = 8'h00;
RAM[16'h2DF7] = 8'h00;
RAM[16'h2DF8] = 8'h00;
RAM[16'h2DF9] = 8'h00;
RAM[16'h2DFA] = 8'h00;
RAM[16'h2DFB] = 8'h00;
RAM[16'h2DFC] = 8'h00;
RAM[16'h2DFD] = 8'h00;
RAM[16'h2DFE] = 8'h00;
RAM[16'h2DFF] = 8'h00;
RAM[16'h2E00] = 8'h00;
RAM[16'h2E01] = 8'h00;
RAM[16'h2E02] = 8'h00;
RAM[16'h2E03] = 8'h00;
RAM[16'h2E04] = 8'h00;
RAM[16'h2E05] = 8'h00;
RAM[16'h2E06] = 8'h00;
RAM[16'h2E07] = 8'h00;
RAM[16'h2E08] = 8'h00;
RAM[16'h2E09] = 8'h00;
RAM[16'h2E0A] = 8'h00;
RAM[16'h2E0B] = 8'h00;
RAM[16'h2E0C] = 8'h00;
RAM[16'h2E0D] = 8'h00;
RAM[16'h2E0E] = 8'h00;
RAM[16'h2E0F] = 8'h00;
RAM[16'h2E10] = 8'h00;
RAM[16'h2E11] = 8'h00;
RAM[16'h2E12] = 8'h00;
RAM[16'h2E13] = 8'h00;
RAM[16'h2E14] = 8'h00;
RAM[16'h2E15] = 8'h00;
RAM[16'h2E16] = 8'h00;
RAM[16'h2E17] = 8'h00;
RAM[16'h2E18] = 8'h00;
RAM[16'h2E19] = 8'h00;
RAM[16'h2E1A] = 8'h00;
RAM[16'h2E1B] = 8'h00;
RAM[16'h2E1C] = 8'h00;
RAM[16'h2E1D] = 8'h00;
RAM[16'h2E1E] = 8'h00;
RAM[16'h2E1F] = 8'h00;
RAM[16'h2E20] = 8'h00;
RAM[16'h2E21] = 8'h00;
RAM[16'h2E22] = 8'h00;
RAM[16'h2E23] = 8'h00;
RAM[16'h2E24] = 8'h00;
RAM[16'h2E25] = 8'h00;
RAM[16'h2E26] = 8'h00;
RAM[16'h2E27] = 8'h00;
RAM[16'h2E28] = 8'h00;
RAM[16'h2E29] = 8'h00;
RAM[16'h2E2A] = 8'h00;
RAM[16'h2E2B] = 8'h00;
RAM[16'h2E2C] = 8'h00;
RAM[16'h2E2D] = 8'h00;
RAM[16'h2E2E] = 8'h00;
RAM[16'h2E2F] = 8'h00;
RAM[16'h2E30] = 8'h00;
RAM[16'h2E31] = 8'h00;
RAM[16'h2E32] = 8'h00;
RAM[16'h2E33] = 8'h00;
RAM[16'h2E34] = 8'h00;
RAM[16'h2E35] = 8'h00;
RAM[16'h2E36] = 8'h00;
RAM[16'h2E37] = 8'h00;
RAM[16'h2E38] = 8'h00;
RAM[16'h2E39] = 8'h00;
RAM[16'h2E3A] = 8'h00;
RAM[16'h2E3B] = 8'h00;
RAM[16'h2E3C] = 8'h00;
RAM[16'h2E3D] = 8'h00;
RAM[16'h2E3E] = 8'h00;
RAM[16'h2E3F] = 8'h00;
RAM[16'h2E40] = 8'h00;
RAM[16'h2E41] = 8'h00;
RAM[16'h2E42] = 8'h00;
RAM[16'h2E43] = 8'h00;
RAM[16'h2E44] = 8'h00;
RAM[16'h2E45] = 8'h00;
RAM[16'h2E46] = 8'h00;
RAM[16'h2E47] = 8'h00;
RAM[16'h2E48] = 8'h00;
RAM[16'h2E49] = 8'h00;
RAM[16'h2E4A] = 8'h00;
RAM[16'h2E4B] = 8'h00;
RAM[16'h2E4C] = 8'h00;
RAM[16'h2E4D] = 8'h00;
RAM[16'h2E4E] = 8'h00;
RAM[16'h2E4F] = 8'h00;
RAM[16'h2E50] = 8'h00;
RAM[16'h2E51] = 8'h00;
RAM[16'h2E52] = 8'h00;
RAM[16'h2E53] = 8'h00;
RAM[16'h2E54] = 8'h00;
RAM[16'h2E55] = 8'h00;
RAM[16'h2E56] = 8'h00;
RAM[16'h2E57] = 8'h00;
RAM[16'h2E58] = 8'h00;
RAM[16'h2E59] = 8'h00;
RAM[16'h2E5A] = 8'h00;
RAM[16'h2E5B] = 8'h00;
RAM[16'h2E5C] = 8'h00;
RAM[16'h2E5D] = 8'h00;
RAM[16'h2E5E] = 8'h00;
RAM[16'h2E5F] = 8'h00;
RAM[16'h2E60] = 8'h00;
RAM[16'h2E61] = 8'h00;
RAM[16'h2E62] = 8'h00;
RAM[16'h2E63] = 8'h00;
RAM[16'h2E64] = 8'h00;
RAM[16'h2E65] = 8'h00;
RAM[16'h2E66] = 8'h00;
RAM[16'h2E67] = 8'h00;
RAM[16'h2E68] = 8'h00;
RAM[16'h2E69] = 8'h00;
RAM[16'h2E6A] = 8'h00;
RAM[16'h2E6B] = 8'h00;
RAM[16'h2E6C] = 8'h00;
RAM[16'h2E6D] = 8'h00;
RAM[16'h2E6E] = 8'h00;
RAM[16'h2E6F] = 8'h00;
RAM[16'h2E70] = 8'h00;
RAM[16'h2E71] = 8'h00;
RAM[16'h2E72] = 8'h00;
RAM[16'h2E73] = 8'h00;
RAM[16'h2E74] = 8'h00;
RAM[16'h2E75] = 8'h00;
RAM[16'h2E76] = 8'h00;
RAM[16'h2E77] = 8'h00;
RAM[16'h2E78] = 8'h00;
RAM[16'h2E79] = 8'h00;
RAM[16'h2E7A] = 8'h00;
RAM[16'h2E7B] = 8'h00;
RAM[16'h2E7C] = 8'h00;
RAM[16'h2E7D] = 8'h00;
RAM[16'h2E7E] = 8'h00;
RAM[16'h2E7F] = 8'h00;
RAM[16'h2E80] = 8'h00;
RAM[16'h2E81] = 8'h00;
RAM[16'h2E82] = 8'h00;
RAM[16'h2E83] = 8'h00;
RAM[16'h2E84] = 8'h00;
RAM[16'h2E85] = 8'h00;
RAM[16'h2E86] = 8'h00;
RAM[16'h2E87] = 8'h00;
RAM[16'h2E88] = 8'h00;
RAM[16'h2E89] = 8'h00;
RAM[16'h2E8A] = 8'h00;
RAM[16'h2E8B] = 8'h00;
RAM[16'h2E8C] = 8'h00;
RAM[16'h2E8D] = 8'h00;
RAM[16'h2E8E] = 8'h00;
RAM[16'h2E8F] = 8'h00;
RAM[16'h2E90] = 8'h00;
RAM[16'h2E91] = 8'h00;
RAM[16'h2E92] = 8'h00;
RAM[16'h2E93] = 8'h00;
RAM[16'h2E94] = 8'h00;
RAM[16'h2E95] = 8'h00;
RAM[16'h2E96] = 8'h00;
RAM[16'h2E97] = 8'h00;
RAM[16'h2E98] = 8'h00;
RAM[16'h2E99] = 8'h00;
RAM[16'h2E9A] = 8'h00;
RAM[16'h2E9B] = 8'h00;
RAM[16'h2E9C] = 8'h00;
RAM[16'h2E9D] = 8'h00;
RAM[16'h2E9E] = 8'h00;
RAM[16'h2E9F] = 8'h00;
RAM[16'h2EA0] = 8'h00;
RAM[16'h2EA1] = 8'h00;
RAM[16'h2EA2] = 8'h00;
RAM[16'h2EA3] = 8'h00;
RAM[16'h2EA4] = 8'h00;
RAM[16'h2EA5] = 8'h00;
RAM[16'h2EA6] = 8'h00;
RAM[16'h2EA7] = 8'h00;
RAM[16'h2EA8] = 8'h00;
RAM[16'h2EA9] = 8'h00;
RAM[16'h2EAA] = 8'h00;
RAM[16'h2EAB] = 8'h00;
RAM[16'h2EAC] = 8'h00;
RAM[16'h2EAD] = 8'h00;
RAM[16'h2EAE] = 8'h00;
RAM[16'h2EAF] = 8'h00;
RAM[16'h2EB0] = 8'h00;
RAM[16'h2EB1] = 8'h00;
RAM[16'h2EB2] = 8'h00;
RAM[16'h2EB3] = 8'h00;
RAM[16'h2EB4] = 8'h00;
RAM[16'h2EB5] = 8'h00;
RAM[16'h2EB6] = 8'h00;
RAM[16'h2EB7] = 8'h00;
RAM[16'h2EB8] = 8'h00;
RAM[16'h2EB9] = 8'h00;
RAM[16'h2EBA] = 8'h00;
RAM[16'h2EBB] = 8'h00;
RAM[16'h2EBC] = 8'h00;
RAM[16'h2EBD] = 8'h00;
RAM[16'h2EBE] = 8'h00;
RAM[16'h2EBF] = 8'h00;
RAM[16'h2EC0] = 8'h00;
RAM[16'h2EC1] = 8'h00;
RAM[16'h2EC2] = 8'h00;
RAM[16'h2EC3] = 8'h00;
RAM[16'h2EC4] = 8'h00;
RAM[16'h2EC5] = 8'h00;
RAM[16'h2EC6] = 8'h00;
RAM[16'h2EC7] = 8'h00;
RAM[16'h2EC8] = 8'h00;
RAM[16'h2EC9] = 8'h00;
RAM[16'h2ECA] = 8'h00;
RAM[16'h2ECB] = 8'h00;
RAM[16'h2ECC] = 8'h00;
RAM[16'h2ECD] = 8'h00;
RAM[16'h2ECE] = 8'h00;
RAM[16'h2ECF] = 8'h00;
RAM[16'h2ED0] = 8'h00;
RAM[16'h2ED1] = 8'h00;
RAM[16'h2ED2] = 8'h00;
RAM[16'h2ED3] = 8'h00;
RAM[16'h2ED4] = 8'h00;
RAM[16'h2ED5] = 8'h00;
RAM[16'h2ED6] = 8'h00;
RAM[16'h2ED7] = 8'h00;
RAM[16'h2ED8] = 8'h00;
RAM[16'h2ED9] = 8'h00;
RAM[16'h2EDA] = 8'h00;
RAM[16'h2EDB] = 8'h00;
RAM[16'h2EDC] = 8'h00;
RAM[16'h2EDD] = 8'h00;
RAM[16'h2EDE] = 8'h00;
RAM[16'h2EDF] = 8'h00;
RAM[16'h2EE0] = 8'h00;
RAM[16'h2EE1] = 8'h00;
RAM[16'h2EE2] = 8'h00;
RAM[16'h2EE3] = 8'h00;
RAM[16'h2EE4] = 8'h00;
RAM[16'h2EE5] = 8'h00;
RAM[16'h2EE6] = 8'h00;
RAM[16'h2EE7] = 8'h00;
RAM[16'h2EE8] = 8'h00;
RAM[16'h2EE9] = 8'h00;
RAM[16'h2EEA] = 8'h00;
RAM[16'h2EEB] = 8'h00;
RAM[16'h2EEC] = 8'h00;
RAM[16'h2EED] = 8'h00;
RAM[16'h2EEE] = 8'h00;
RAM[16'h2EEF] = 8'h00;
RAM[16'h2EF0] = 8'h00;
RAM[16'h2EF1] = 8'h00;
RAM[16'h2EF2] = 8'h00;
RAM[16'h2EF3] = 8'h00;
RAM[16'h2EF4] = 8'h00;
RAM[16'h2EF5] = 8'h00;
RAM[16'h2EF6] = 8'h00;
RAM[16'h2EF7] = 8'h00;
RAM[16'h2EF8] = 8'h00;
RAM[16'h2EF9] = 8'h00;
RAM[16'h2EFA] = 8'h00;
RAM[16'h2EFB] = 8'h00;
RAM[16'h2EFC] = 8'h00;
RAM[16'h2EFD] = 8'h00;
RAM[16'h2EFE] = 8'h00;
RAM[16'h2EFF] = 8'h00;
RAM[16'h2F00] = 8'h00;
RAM[16'h2F01] = 8'h00;
RAM[16'h2F02] = 8'h00;
RAM[16'h2F03] = 8'h00;
RAM[16'h2F04] = 8'h00;
RAM[16'h2F05] = 8'h00;
RAM[16'h2F06] = 8'h00;
RAM[16'h2F07] = 8'h00;
RAM[16'h2F08] = 8'h00;
RAM[16'h2F09] = 8'h00;
RAM[16'h2F0A] = 8'h00;
RAM[16'h2F0B] = 8'h00;
RAM[16'h2F0C] = 8'h00;
RAM[16'h2F0D] = 8'h00;
RAM[16'h2F0E] = 8'h00;
RAM[16'h2F0F] = 8'h00;
RAM[16'h2F10] = 8'h00;
RAM[16'h2F11] = 8'h00;
RAM[16'h2F12] = 8'h00;
RAM[16'h2F13] = 8'h00;
RAM[16'h2F14] = 8'h00;
RAM[16'h2F15] = 8'h00;
RAM[16'h2F16] = 8'h00;
RAM[16'h2F17] = 8'h00;
RAM[16'h2F18] = 8'h00;
RAM[16'h2F19] = 8'h00;
RAM[16'h2F1A] = 8'h00;
RAM[16'h2F1B] = 8'h00;
RAM[16'h2F1C] = 8'h00;
RAM[16'h2F1D] = 8'h00;
RAM[16'h2F1E] = 8'h00;
RAM[16'h2F1F] = 8'h00;
RAM[16'h2F20] = 8'h00;
RAM[16'h2F21] = 8'h00;
RAM[16'h2F22] = 8'h00;
RAM[16'h2F23] = 8'h00;
RAM[16'h2F24] = 8'h00;
RAM[16'h2F25] = 8'h00;
RAM[16'h2F26] = 8'h00;
RAM[16'h2F27] = 8'h00;
RAM[16'h2F28] = 8'h00;
RAM[16'h2F29] = 8'h00;
RAM[16'h2F2A] = 8'h00;
RAM[16'h2F2B] = 8'h00;
RAM[16'h2F2C] = 8'h00;
RAM[16'h2F2D] = 8'h00;
RAM[16'h2F2E] = 8'h00;
RAM[16'h2F2F] = 8'h00;
RAM[16'h2F30] = 8'h00;
RAM[16'h2F31] = 8'h00;
RAM[16'h2F32] = 8'h00;
RAM[16'h2F33] = 8'h00;
RAM[16'h2F34] = 8'h00;
RAM[16'h2F35] = 8'h00;
RAM[16'h2F36] = 8'h00;
RAM[16'h2F37] = 8'h00;
RAM[16'h2F38] = 8'h00;
RAM[16'h2F39] = 8'h00;
RAM[16'h2F3A] = 8'h00;
RAM[16'h2F3B] = 8'h00;
RAM[16'h2F3C] = 8'h00;
RAM[16'h2F3D] = 8'h00;
RAM[16'h2F3E] = 8'h00;
RAM[16'h2F3F] = 8'h00;
RAM[16'h2F40] = 8'h00;
RAM[16'h2F41] = 8'h00;
RAM[16'h2F42] = 8'h00;
RAM[16'h2F43] = 8'h00;
RAM[16'h2F44] = 8'h00;
RAM[16'h2F45] = 8'h00;
RAM[16'h2F46] = 8'h00;
RAM[16'h2F47] = 8'h00;
RAM[16'h2F48] = 8'h00;
RAM[16'h2F49] = 8'h00;
RAM[16'h2F4A] = 8'h00;
RAM[16'h2F4B] = 8'h00;
RAM[16'h2F4C] = 8'h00;
RAM[16'h2F4D] = 8'h00;
RAM[16'h2F4E] = 8'h00;
RAM[16'h2F4F] = 8'h00;
RAM[16'h2F50] = 8'h00;
RAM[16'h2F51] = 8'h00;
RAM[16'h2F52] = 8'h00;
RAM[16'h2F53] = 8'h00;
RAM[16'h2F54] = 8'h00;
RAM[16'h2F55] = 8'h00;
RAM[16'h2F56] = 8'h00;
RAM[16'h2F57] = 8'h00;
RAM[16'h2F58] = 8'h00;
RAM[16'h2F59] = 8'h00;
RAM[16'h2F5A] = 8'h00;
RAM[16'h2F5B] = 8'h00;
RAM[16'h2F5C] = 8'h00;
RAM[16'h2F5D] = 8'h00;
RAM[16'h2F5E] = 8'h00;
RAM[16'h2F5F] = 8'h00;
RAM[16'h2F60] = 8'h00;
RAM[16'h2F61] = 8'h00;
RAM[16'h2F62] = 8'h00;
RAM[16'h2F63] = 8'h00;
RAM[16'h2F64] = 8'h00;
RAM[16'h2F65] = 8'h00;
RAM[16'h2F66] = 8'h00;
RAM[16'h2F67] = 8'h00;
RAM[16'h2F68] = 8'h00;
RAM[16'h2F69] = 8'h00;
RAM[16'h2F6A] = 8'h00;
RAM[16'h2F6B] = 8'h00;
RAM[16'h2F6C] = 8'h00;
RAM[16'h2F6D] = 8'h00;
RAM[16'h2F6E] = 8'h00;
RAM[16'h2F6F] = 8'h00;
RAM[16'h2F70] = 8'h00;
RAM[16'h2F71] = 8'h00;
RAM[16'h2F72] = 8'h00;
RAM[16'h2F73] = 8'h00;
RAM[16'h2F74] = 8'h00;
RAM[16'h2F75] = 8'h00;
RAM[16'h2F76] = 8'h00;
RAM[16'h2F77] = 8'h00;
RAM[16'h2F78] = 8'h00;
RAM[16'h2F79] = 8'h00;
RAM[16'h2F7A] = 8'h00;
RAM[16'h2F7B] = 8'h00;
RAM[16'h2F7C] = 8'h00;
RAM[16'h2F7D] = 8'h00;
RAM[16'h2F7E] = 8'h00;
RAM[16'h2F7F] = 8'h00;
RAM[16'h2F80] = 8'h00;
RAM[16'h2F81] = 8'h00;
RAM[16'h2F82] = 8'h00;
RAM[16'h2F83] = 8'h00;
RAM[16'h2F84] = 8'h00;
RAM[16'h2F85] = 8'h00;
RAM[16'h2F86] = 8'h00;
RAM[16'h2F87] = 8'h00;
RAM[16'h2F88] = 8'h00;
RAM[16'h2F89] = 8'h00;
RAM[16'h2F8A] = 8'h00;
RAM[16'h2F8B] = 8'h00;
RAM[16'h2F8C] = 8'h00;
RAM[16'h2F8D] = 8'h00;
RAM[16'h2F8E] = 8'h00;
RAM[16'h2F8F] = 8'h00;
RAM[16'h2F90] = 8'h00;
RAM[16'h2F91] = 8'h00;
RAM[16'h2F92] = 8'h00;
RAM[16'h2F93] = 8'h00;
RAM[16'h2F94] = 8'h00;
RAM[16'h2F95] = 8'h00;
RAM[16'h2F96] = 8'h00;
RAM[16'h2F97] = 8'h00;
RAM[16'h2F98] = 8'h00;
RAM[16'h2F99] = 8'h00;
RAM[16'h2F9A] = 8'h00;
RAM[16'h2F9B] = 8'h00;
RAM[16'h2F9C] = 8'h00;
RAM[16'h2F9D] = 8'h00;
RAM[16'h2F9E] = 8'h00;
RAM[16'h2F9F] = 8'h00;
RAM[16'h2FA0] = 8'h00;
RAM[16'h2FA1] = 8'h00;
RAM[16'h2FA2] = 8'h00;
RAM[16'h2FA3] = 8'h00;
RAM[16'h2FA4] = 8'h00;
RAM[16'h2FA5] = 8'h00;
RAM[16'h2FA6] = 8'h00;
RAM[16'h2FA7] = 8'h00;
RAM[16'h2FA8] = 8'h00;
RAM[16'h2FA9] = 8'h00;
RAM[16'h2FAA] = 8'h00;
RAM[16'h2FAB] = 8'h00;
RAM[16'h2FAC] = 8'h00;
RAM[16'h2FAD] = 8'h00;
RAM[16'h2FAE] = 8'h00;
RAM[16'h2FAF] = 8'h00;
RAM[16'h2FB0] = 8'h00;
RAM[16'h2FB1] = 8'h00;
RAM[16'h2FB2] = 8'h00;
RAM[16'h2FB3] = 8'h00;
RAM[16'h2FB4] = 8'h00;
RAM[16'h2FB5] = 8'h00;
RAM[16'h2FB6] = 8'h00;
RAM[16'h2FB7] = 8'h00;
RAM[16'h2FB8] = 8'h00;
RAM[16'h2FB9] = 8'h00;
RAM[16'h2FBA] = 8'h00;
RAM[16'h2FBB] = 8'h00;
RAM[16'h2FBC] = 8'h00;
RAM[16'h2FBD] = 8'h00;
RAM[16'h2FBE] = 8'h00;
RAM[16'h2FBF] = 8'h00;
RAM[16'h2FC0] = 8'h00;
RAM[16'h2FC1] = 8'h00;
RAM[16'h2FC2] = 8'h00;
RAM[16'h2FC3] = 8'h00;
RAM[16'h2FC4] = 8'h00;
RAM[16'h2FC5] = 8'h00;
RAM[16'h2FC6] = 8'h00;
RAM[16'h2FC7] = 8'h00;
RAM[16'h2FC8] = 8'h00;
RAM[16'h2FC9] = 8'h00;
RAM[16'h2FCA] = 8'h00;
RAM[16'h2FCB] = 8'h00;
RAM[16'h2FCC] = 8'h00;
RAM[16'h2FCD] = 8'h00;
RAM[16'h2FCE] = 8'h00;
RAM[16'h2FCF] = 8'h00;
RAM[16'h2FD0] = 8'h00;
RAM[16'h2FD1] = 8'h00;
RAM[16'h2FD2] = 8'h00;
RAM[16'h2FD3] = 8'h00;
RAM[16'h2FD4] = 8'h00;
RAM[16'h2FD5] = 8'h00;
RAM[16'h2FD6] = 8'h00;
RAM[16'h2FD7] = 8'h00;
RAM[16'h2FD8] = 8'h00;
RAM[16'h2FD9] = 8'h00;
RAM[16'h2FDA] = 8'h00;
RAM[16'h2FDB] = 8'h00;
RAM[16'h2FDC] = 8'h00;
RAM[16'h2FDD] = 8'h00;
RAM[16'h2FDE] = 8'h00;
RAM[16'h2FDF] = 8'h00;
RAM[16'h2FE0] = 8'h00;
RAM[16'h2FE1] = 8'h00;
RAM[16'h2FE2] = 8'h00;
RAM[16'h2FE3] = 8'h00;
RAM[16'h2FE4] = 8'h00;
RAM[16'h2FE5] = 8'h00;
RAM[16'h2FE6] = 8'h00;
RAM[16'h2FE7] = 8'h00;
RAM[16'h2FE8] = 8'h00;
RAM[16'h2FE9] = 8'h00;
RAM[16'h2FEA] = 8'h00;
RAM[16'h2FEB] = 8'h00;
RAM[16'h2FEC] = 8'h00;
RAM[16'h2FED] = 8'h00;
RAM[16'h2FEE] = 8'h00;
RAM[16'h2FEF] = 8'h00;
RAM[16'h2FF0] = 8'h00;
RAM[16'h2FF1] = 8'h00;
RAM[16'h2FF2] = 8'h00;
RAM[16'h2FF3] = 8'h00;
RAM[16'h2FF4] = 8'h00;
RAM[16'h2FF5] = 8'h00;
RAM[16'h2FF6] = 8'h00;
RAM[16'h2FF7] = 8'h00;
RAM[16'h2FF8] = 8'h00;
RAM[16'h2FF9] = 8'h00;
RAM[16'h2FFA] = 8'h00;
RAM[16'h2FFB] = 8'h00;
RAM[16'h2FFC] = 8'h00;
RAM[16'h2FFD] = 8'h00;
RAM[16'h2FFE] = 8'h00;
RAM[16'h2FFF] = 8'h00;
RAM[16'h3000] = 8'h00;
RAM[16'h3001] = 8'h00;
RAM[16'h3002] = 8'h00;
RAM[16'h3003] = 8'h00;
RAM[16'h3004] = 8'h00;
RAM[16'h3005] = 8'h00;
RAM[16'h3006] = 8'h00;
RAM[16'h3007] = 8'h00;
RAM[16'h3008] = 8'h00;
RAM[16'h3009] = 8'h00;
RAM[16'h300A] = 8'h00;
RAM[16'h300B] = 8'h00;
RAM[16'h300C] = 8'h00;
RAM[16'h300D] = 8'h00;
RAM[16'h300E] = 8'h00;
RAM[16'h300F] = 8'h00;
RAM[16'h3010] = 8'h00;
RAM[16'h3011] = 8'h00;
RAM[16'h3012] = 8'h00;
RAM[16'h3013] = 8'h00;
RAM[16'h3014] = 8'h00;
RAM[16'h3015] = 8'h00;
RAM[16'h3016] = 8'h00;
RAM[16'h3017] = 8'h00;
RAM[16'h3018] = 8'h00;
RAM[16'h3019] = 8'h00;
RAM[16'h301A] = 8'h00;
RAM[16'h301B] = 8'h00;
RAM[16'h301C] = 8'h00;
RAM[16'h301D] = 8'h00;
RAM[16'h301E] = 8'h00;
RAM[16'h301F] = 8'h00;
RAM[16'h3020] = 8'h00;
RAM[16'h3021] = 8'h00;
RAM[16'h3022] = 8'h00;
RAM[16'h3023] = 8'h00;
RAM[16'h3024] = 8'h00;
RAM[16'h3025] = 8'h00;
RAM[16'h3026] = 8'h00;
RAM[16'h3027] = 8'h00;
RAM[16'h3028] = 8'h00;
RAM[16'h3029] = 8'h00;
RAM[16'h302A] = 8'h00;
RAM[16'h302B] = 8'h00;
RAM[16'h302C] = 8'h00;
RAM[16'h302D] = 8'h00;
RAM[16'h302E] = 8'h00;
RAM[16'h302F] = 8'h00;
RAM[16'h3030] = 8'h00;
RAM[16'h3031] = 8'h00;
RAM[16'h3032] = 8'h00;
RAM[16'h3033] = 8'h00;
RAM[16'h3034] = 8'h00;
RAM[16'h3035] = 8'h00;
RAM[16'h3036] = 8'h00;
RAM[16'h3037] = 8'h00;
RAM[16'h3038] = 8'h00;
RAM[16'h3039] = 8'h00;
RAM[16'h303A] = 8'h00;
RAM[16'h303B] = 8'h00;
RAM[16'h303C] = 8'h00;
RAM[16'h303D] = 8'h00;
RAM[16'h303E] = 8'h00;
RAM[16'h303F] = 8'h00;
RAM[16'h3040] = 8'h00;
RAM[16'h3041] = 8'h00;
RAM[16'h3042] = 8'h00;
RAM[16'h3043] = 8'h00;
RAM[16'h3044] = 8'h00;
RAM[16'h3045] = 8'h00;
RAM[16'h3046] = 8'h00;
RAM[16'h3047] = 8'h00;
RAM[16'h3048] = 8'h00;
RAM[16'h3049] = 8'h00;
RAM[16'h304A] = 8'h00;
RAM[16'h304B] = 8'h00;
RAM[16'h304C] = 8'h00;
RAM[16'h304D] = 8'h00;
RAM[16'h304E] = 8'h00;
RAM[16'h304F] = 8'h00;
RAM[16'h3050] = 8'h00;
RAM[16'h3051] = 8'h00;
RAM[16'h3052] = 8'h00;
RAM[16'h3053] = 8'h00;
RAM[16'h3054] = 8'h00;
RAM[16'h3055] = 8'h00;
RAM[16'h3056] = 8'h00;
RAM[16'h3057] = 8'h00;
RAM[16'h3058] = 8'h00;
RAM[16'h3059] = 8'h00;
RAM[16'h305A] = 8'h00;
RAM[16'h305B] = 8'h00;
RAM[16'h305C] = 8'h00;
RAM[16'h305D] = 8'h00;
RAM[16'h305E] = 8'h00;
RAM[16'h305F] = 8'h00;
RAM[16'h3060] = 8'h00;
RAM[16'h3061] = 8'h00;
RAM[16'h3062] = 8'h00;
RAM[16'h3063] = 8'h00;
RAM[16'h3064] = 8'h00;
RAM[16'h3065] = 8'h00;
RAM[16'h3066] = 8'h00;
RAM[16'h3067] = 8'h00;
RAM[16'h3068] = 8'h00;
RAM[16'h3069] = 8'h00;
RAM[16'h306A] = 8'h00;
RAM[16'h306B] = 8'h00;
RAM[16'h306C] = 8'h00;
RAM[16'h306D] = 8'h00;
RAM[16'h306E] = 8'h00;
RAM[16'h306F] = 8'h00;
RAM[16'h3070] = 8'h00;
RAM[16'h3071] = 8'h00;
RAM[16'h3072] = 8'h00;
RAM[16'h3073] = 8'h00;
RAM[16'h3074] = 8'h00;
RAM[16'h3075] = 8'h00;
RAM[16'h3076] = 8'h00;
RAM[16'h3077] = 8'h00;
RAM[16'h3078] = 8'h00;
RAM[16'h3079] = 8'h00;
RAM[16'h307A] = 8'h00;
RAM[16'h307B] = 8'h00;
RAM[16'h307C] = 8'h00;
RAM[16'h307D] = 8'h00;
RAM[16'h307E] = 8'h00;
RAM[16'h307F] = 8'h00;
RAM[16'h3080] = 8'h00;
RAM[16'h3081] = 8'h00;
RAM[16'h3082] = 8'h00;
RAM[16'h3083] = 8'h00;
RAM[16'h3084] = 8'h00;
RAM[16'h3085] = 8'h00;
RAM[16'h3086] = 8'h00;
RAM[16'h3087] = 8'h00;
RAM[16'h3088] = 8'h00;
RAM[16'h3089] = 8'h00;
RAM[16'h308A] = 8'h00;
RAM[16'h308B] = 8'h00;
RAM[16'h308C] = 8'h00;
RAM[16'h308D] = 8'h00;
RAM[16'h308E] = 8'h00;
RAM[16'h308F] = 8'h00;
RAM[16'h3090] = 8'h00;
RAM[16'h3091] = 8'h00;
RAM[16'h3092] = 8'h00;
RAM[16'h3093] = 8'h00;
RAM[16'h3094] = 8'h00;
RAM[16'h3095] = 8'h00;
RAM[16'h3096] = 8'h00;
RAM[16'h3097] = 8'h00;
RAM[16'h3098] = 8'h00;
RAM[16'h3099] = 8'h00;
RAM[16'h309A] = 8'h00;
RAM[16'h309B] = 8'h00;
RAM[16'h309C] = 8'h00;
RAM[16'h309D] = 8'h00;
RAM[16'h309E] = 8'h00;
RAM[16'h309F] = 8'h00;
RAM[16'h30A0] = 8'h00;
RAM[16'h30A1] = 8'h00;
RAM[16'h30A2] = 8'h00;
RAM[16'h30A3] = 8'h00;
RAM[16'h30A4] = 8'h00;
RAM[16'h30A5] = 8'h00;
RAM[16'h30A6] = 8'h00;
RAM[16'h30A7] = 8'h00;
RAM[16'h30A8] = 8'h00;
RAM[16'h30A9] = 8'h00;
RAM[16'h30AA] = 8'h00;
RAM[16'h30AB] = 8'h00;
RAM[16'h30AC] = 8'h00;
RAM[16'h30AD] = 8'h00;
RAM[16'h30AE] = 8'h00;
RAM[16'h30AF] = 8'h00;
RAM[16'h30B0] = 8'h00;
RAM[16'h30B1] = 8'h00;
RAM[16'h30B2] = 8'h00;
RAM[16'h30B3] = 8'h00;
RAM[16'h30B4] = 8'h00;
RAM[16'h30B5] = 8'h00;
RAM[16'h30B6] = 8'h00;
RAM[16'h30B7] = 8'h00;
RAM[16'h30B8] = 8'h00;
RAM[16'h30B9] = 8'h00;
RAM[16'h30BA] = 8'h00;
RAM[16'h30BB] = 8'h00;
RAM[16'h30BC] = 8'h00;
RAM[16'h30BD] = 8'h00;
RAM[16'h30BE] = 8'h00;
RAM[16'h30BF] = 8'h00;
RAM[16'h30C0] = 8'h00;
RAM[16'h30C1] = 8'h00;
RAM[16'h30C2] = 8'h00;
RAM[16'h30C3] = 8'h00;
RAM[16'h30C4] = 8'h00;
RAM[16'h30C5] = 8'h00;
RAM[16'h30C6] = 8'h00;
RAM[16'h30C7] = 8'h00;
RAM[16'h30C8] = 8'h00;
RAM[16'h30C9] = 8'h00;
RAM[16'h30CA] = 8'h00;
RAM[16'h30CB] = 8'h00;
RAM[16'h30CC] = 8'h00;
RAM[16'h30CD] = 8'h00;
RAM[16'h30CE] = 8'h00;
RAM[16'h30CF] = 8'h00;
RAM[16'h30D0] = 8'h00;
RAM[16'h30D1] = 8'h00;
RAM[16'h30D2] = 8'h00;
RAM[16'h30D3] = 8'h00;
RAM[16'h30D4] = 8'h00;
RAM[16'h30D5] = 8'h00;
RAM[16'h30D6] = 8'h00;
RAM[16'h30D7] = 8'h00;
RAM[16'h30D8] = 8'h00;
RAM[16'h30D9] = 8'h00;
RAM[16'h30DA] = 8'h00;
RAM[16'h30DB] = 8'h00;
RAM[16'h30DC] = 8'h00;
RAM[16'h30DD] = 8'h00;
RAM[16'h30DE] = 8'h00;
RAM[16'h30DF] = 8'h00;
RAM[16'h30E0] = 8'h00;
RAM[16'h30E1] = 8'h00;
RAM[16'h30E2] = 8'h00;
RAM[16'h30E3] = 8'h00;
RAM[16'h30E4] = 8'h00;
RAM[16'h30E5] = 8'h00;
RAM[16'h30E6] = 8'h00;
RAM[16'h30E7] = 8'h00;
RAM[16'h30E8] = 8'h00;
RAM[16'h30E9] = 8'h00;
RAM[16'h30EA] = 8'h00;
RAM[16'h30EB] = 8'h00;
RAM[16'h30EC] = 8'h00;
RAM[16'h30ED] = 8'h00;
RAM[16'h30EE] = 8'h00;
RAM[16'h30EF] = 8'h00;
RAM[16'h30F0] = 8'h00;
RAM[16'h30F1] = 8'h00;
RAM[16'h30F2] = 8'h00;
RAM[16'h30F3] = 8'h00;
RAM[16'h30F4] = 8'h00;
RAM[16'h30F5] = 8'h00;
RAM[16'h30F6] = 8'h00;
RAM[16'h30F7] = 8'h00;
RAM[16'h30F8] = 8'h00;
RAM[16'h30F9] = 8'h00;
RAM[16'h30FA] = 8'h00;
RAM[16'h30FB] = 8'h00;
RAM[16'h30FC] = 8'h00;
RAM[16'h30FD] = 8'h00;
RAM[16'h30FE] = 8'h00;
RAM[16'h30FF] = 8'h00;
RAM[16'h3100] = 8'h00;
RAM[16'h3101] = 8'h00;
RAM[16'h3102] = 8'h00;
RAM[16'h3103] = 8'h00;
RAM[16'h3104] = 8'h00;
RAM[16'h3105] = 8'h00;
RAM[16'h3106] = 8'h00;
RAM[16'h3107] = 8'h00;
RAM[16'h3108] = 8'h00;
RAM[16'h3109] = 8'h00;
RAM[16'h310A] = 8'h00;
RAM[16'h310B] = 8'h00;
RAM[16'h310C] = 8'h00;
RAM[16'h310D] = 8'h00;
RAM[16'h310E] = 8'h00;
RAM[16'h310F] = 8'h00;
RAM[16'h3110] = 8'h00;
RAM[16'h3111] = 8'h00;
RAM[16'h3112] = 8'h00;
RAM[16'h3113] = 8'h00;
RAM[16'h3114] = 8'h00;
RAM[16'h3115] = 8'h00;
RAM[16'h3116] = 8'h00;
RAM[16'h3117] = 8'h00;
RAM[16'h3118] = 8'h00;
RAM[16'h3119] = 8'h00;
RAM[16'h311A] = 8'h00;
RAM[16'h311B] = 8'h00;
RAM[16'h311C] = 8'h00;
RAM[16'h311D] = 8'h00;
RAM[16'h311E] = 8'h00;
RAM[16'h311F] = 8'h00;
RAM[16'h3120] = 8'h00;
RAM[16'h3121] = 8'h00;
RAM[16'h3122] = 8'h00;
RAM[16'h3123] = 8'h00;
RAM[16'h3124] = 8'h00;
RAM[16'h3125] = 8'h00;
RAM[16'h3126] = 8'h00;
RAM[16'h3127] = 8'h00;
RAM[16'h3128] = 8'h00;
RAM[16'h3129] = 8'h00;
RAM[16'h312A] = 8'h00;
RAM[16'h312B] = 8'h00;
RAM[16'h312C] = 8'h00;
RAM[16'h312D] = 8'h00;
RAM[16'h312E] = 8'h00;
RAM[16'h312F] = 8'h00;
RAM[16'h3130] = 8'h00;
RAM[16'h3131] = 8'h00;
RAM[16'h3132] = 8'h00;
RAM[16'h3133] = 8'h00;
RAM[16'h3134] = 8'h00;
RAM[16'h3135] = 8'h00;
RAM[16'h3136] = 8'h00;
RAM[16'h3137] = 8'h00;
RAM[16'h3138] = 8'h00;
RAM[16'h3139] = 8'h00;
RAM[16'h313A] = 8'h00;
RAM[16'h313B] = 8'h00;
RAM[16'h313C] = 8'h00;
RAM[16'h313D] = 8'h00;
RAM[16'h313E] = 8'h00;
RAM[16'h313F] = 8'h00;
RAM[16'h3140] = 8'h00;
RAM[16'h3141] = 8'h00;
RAM[16'h3142] = 8'h00;
RAM[16'h3143] = 8'h00;
RAM[16'h3144] = 8'h00;
RAM[16'h3145] = 8'h00;
RAM[16'h3146] = 8'h00;
RAM[16'h3147] = 8'h00;
RAM[16'h3148] = 8'h00;
RAM[16'h3149] = 8'h00;
RAM[16'h314A] = 8'h00;
RAM[16'h314B] = 8'h00;
RAM[16'h314C] = 8'h00;
RAM[16'h314D] = 8'h00;
RAM[16'h314E] = 8'h00;
RAM[16'h314F] = 8'h00;
RAM[16'h3150] = 8'h00;
RAM[16'h3151] = 8'h00;
RAM[16'h3152] = 8'h00;
RAM[16'h3153] = 8'h00;
RAM[16'h3154] = 8'h00;
RAM[16'h3155] = 8'h00;
RAM[16'h3156] = 8'h00;
RAM[16'h3157] = 8'h00;
RAM[16'h3158] = 8'h00;
RAM[16'h3159] = 8'h00;
RAM[16'h315A] = 8'h00;
RAM[16'h315B] = 8'h00;
RAM[16'h315C] = 8'h00;
RAM[16'h315D] = 8'h00;
RAM[16'h315E] = 8'h00;
RAM[16'h315F] = 8'h00;
RAM[16'h3160] = 8'h00;
RAM[16'h3161] = 8'h00;
RAM[16'h3162] = 8'h00;
RAM[16'h3163] = 8'h00;
RAM[16'h3164] = 8'h00;
RAM[16'h3165] = 8'h00;
RAM[16'h3166] = 8'h00;
RAM[16'h3167] = 8'h00;
RAM[16'h3168] = 8'h00;
RAM[16'h3169] = 8'h00;
RAM[16'h316A] = 8'h00;
RAM[16'h316B] = 8'h00;
RAM[16'h316C] = 8'h00;
RAM[16'h316D] = 8'h00;
RAM[16'h316E] = 8'h00;
RAM[16'h316F] = 8'h00;
RAM[16'h3170] = 8'h00;
RAM[16'h3171] = 8'h00;
RAM[16'h3172] = 8'h00;
RAM[16'h3173] = 8'h00;
RAM[16'h3174] = 8'h00;
RAM[16'h3175] = 8'h00;
RAM[16'h3176] = 8'h00;
RAM[16'h3177] = 8'h00;
RAM[16'h3178] = 8'h00;
RAM[16'h3179] = 8'h00;
RAM[16'h317A] = 8'h00;
RAM[16'h317B] = 8'h00;
RAM[16'h317C] = 8'h00;
RAM[16'h317D] = 8'h00;
RAM[16'h317E] = 8'h00;
RAM[16'h317F] = 8'h00;
RAM[16'h3180] = 8'h00;
RAM[16'h3181] = 8'h00;
RAM[16'h3182] = 8'h00;
RAM[16'h3183] = 8'h00;
RAM[16'h3184] = 8'h00;
RAM[16'h3185] = 8'h00;
RAM[16'h3186] = 8'h00;
RAM[16'h3187] = 8'h00;
RAM[16'h3188] = 8'h00;
RAM[16'h3189] = 8'h00;
RAM[16'h318A] = 8'h00;
RAM[16'h318B] = 8'h00;
RAM[16'h318C] = 8'h00;
RAM[16'h318D] = 8'h00;
RAM[16'h318E] = 8'h00;
RAM[16'h318F] = 8'h00;
RAM[16'h3190] = 8'h00;
RAM[16'h3191] = 8'h00;
RAM[16'h3192] = 8'h00;
RAM[16'h3193] = 8'h00;
RAM[16'h3194] = 8'h00;
RAM[16'h3195] = 8'h00;
RAM[16'h3196] = 8'h00;
RAM[16'h3197] = 8'h00;
RAM[16'h3198] = 8'h00;
RAM[16'h3199] = 8'h00;
RAM[16'h319A] = 8'h00;
RAM[16'h319B] = 8'h00;
RAM[16'h319C] = 8'h00;
RAM[16'h319D] = 8'h00;
RAM[16'h319E] = 8'h00;
RAM[16'h319F] = 8'h00;
RAM[16'h31A0] = 8'h00;
RAM[16'h31A1] = 8'h00;
RAM[16'h31A2] = 8'h00;
RAM[16'h31A3] = 8'h00;
RAM[16'h31A4] = 8'h00;
RAM[16'h31A5] = 8'h00;
RAM[16'h31A6] = 8'h00;
RAM[16'h31A7] = 8'h00;
RAM[16'h31A8] = 8'h00;
RAM[16'h31A9] = 8'h00;
RAM[16'h31AA] = 8'h00;
RAM[16'h31AB] = 8'h00;
RAM[16'h31AC] = 8'h00;
RAM[16'h31AD] = 8'h00;
RAM[16'h31AE] = 8'h00;
RAM[16'h31AF] = 8'h00;
RAM[16'h31B0] = 8'h00;
RAM[16'h31B1] = 8'h00;
RAM[16'h31B2] = 8'h00;
RAM[16'h31B3] = 8'h00;
RAM[16'h31B4] = 8'h00;
RAM[16'h31B5] = 8'h00;
RAM[16'h31B6] = 8'h00;
RAM[16'h31B7] = 8'h00;
RAM[16'h31B8] = 8'h00;
RAM[16'h31B9] = 8'h00;
RAM[16'h31BA] = 8'h00;
RAM[16'h31BB] = 8'h00;
RAM[16'h31BC] = 8'h00;
RAM[16'h31BD] = 8'h00;
RAM[16'h31BE] = 8'h00;
RAM[16'h31BF] = 8'h00;
RAM[16'h31C0] = 8'h00;
RAM[16'h31C1] = 8'h00;
RAM[16'h31C2] = 8'h00;
RAM[16'h31C3] = 8'h00;
RAM[16'h31C4] = 8'h00;
RAM[16'h31C5] = 8'h00;
RAM[16'h31C6] = 8'h00;
RAM[16'h31C7] = 8'h00;
RAM[16'h31C8] = 8'h00;
RAM[16'h31C9] = 8'h00;
RAM[16'h31CA] = 8'h00;
RAM[16'h31CB] = 8'h00;
RAM[16'h31CC] = 8'h00;
RAM[16'h31CD] = 8'h00;
RAM[16'h31CE] = 8'h00;
RAM[16'h31CF] = 8'h00;
RAM[16'h31D0] = 8'h00;
RAM[16'h31D1] = 8'h00;
RAM[16'h31D2] = 8'h00;
RAM[16'h31D3] = 8'h00;
RAM[16'h31D4] = 8'h00;
RAM[16'h31D5] = 8'h00;
RAM[16'h31D6] = 8'h00;
RAM[16'h31D7] = 8'h00;
RAM[16'h31D8] = 8'h00;
RAM[16'h31D9] = 8'h00;
RAM[16'h31DA] = 8'h00;
RAM[16'h31DB] = 8'h00;
RAM[16'h31DC] = 8'h00;
RAM[16'h31DD] = 8'h00;
RAM[16'h31DE] = 8'h00;
RAM[16'h31DF] = 8'h00;
RAM[16'h31E0] = 8'h00;
RAM[16'h31E1] = 8'h00;
RAM[16'h31E2] = 8'h00;
RAM[16'h31E3] = 8'h00;
RAM[16'h31E4] = 8'h00;
RAM[16'h31E5] = 8'h00;
RAM[16'h31E6] = 8'h00;
RAM[16'h31E7] = 8'h00;
RAM[16'h31E8] = 8'h00;
RAM[16'h31E9] = 8'h00;
RAM[16'h31EA] = 8'h00;
RAM[16'h31EB] = 8'h00;
RAM[16'h31EC] = 8'h00;
RAM[16'h31ED] = 8'h00;
RAM[16'h31EE] = 8'h00;
RAM[16'h31EF] = 8'h00;
RAM[16'h31F0] = 8'h00;
RAM[16'h31F1] = 8'h00;
RAM[16'h31F2] = 8'h00;
RAM[16'h31F3] = 8'h00;
RAM[16'h31F4] = 8'h00;
RAM[16'h31F5] = 8'h00;
RAM[16'h31F6] = 8'h00;
RAM[16'h31F7] = 8'h00;
RAM[16'h31F8] = 8'h00;
RAM[16'h31F9] = 8'h00;
RAM[16'h31FA] = 8'h00;
RAM[16'h31FB] = 8'h00;
RAM[16'h31FC] = 8'h00;
RAM[16'h31FD] = 8'h00;
RAM[16'h31FE] = 8'h00;
RAM[16'h31FF] = 8'h00;
RAM[16'h3200] = 8'h00;
RAM[16'h3201] = 8'h00;
RAM[16'h3202] = 8'h00;
RAM[16'h3203] = 8'h00;
RAM[16'h3204] = 8'h00;
RAM[16'h3205] = 8'h00;
RAM[16'h3206] = 8'h00;
RAM[16'h3207] = 8'h00;
RAM[16'h3208] = 8'h00;
RAM[16'h3209] = 8'h00;
RAM[16'h320A] = 8'h00;
RAM[16'h320B] = 8'h00;
RAM[16'h320C] = 8'h00;
RAM[16'h320D] = 8'h00;
RAM[16'h320E] = 8'h00;
RAM[16'h320F] = 8'h00;
RAM[16'h3210] = 8'h00;
RAM[16'h3211] = 8'h00;
RAM[16'h3212] = 8'h00;
RAM[16'h3213] = 8'h00;
RAM[16'h3214] = 8'h00;
RAM[16'h3215] = 8'h00;
RAM[16'h3216] = 8'h00;
RAM[16'h3217] = 8'h00;
RAM[16'h3218] = 8'h00;
RAM[16'h3219] = 8'h00;
RAM[16'h321A] = 8'h00;
RAM[16'h321B] = 8'h00;
RAM[16'h321C] = 8'h00;
RAM[16'h321D] = 8'h00;
RAM[16'h321E] = 8'h00;
RAM[16'h321F] = 8'h00;
RAM[16'h3220] = 8'h00;
RAM[16'h3221] = 8'h00;
RAM[16'h3222] = 8'h00;
RAM[16'h3223] = 8'h00;
RAM[16'h3224] = 8'h00;
RAM[16'h3225] = 8'h00;
RAM[16'h3226] = 8'h00;
RAM[16'h3227] = 8'h00;
RAM[16'h3228] = 8'h00;
RAM[16'h3229] = 8'h00;
RAM[16'h322A] = 8'h00;
RAM[16'h322B] = 8'h00;
RAM[16'h322C] = 8'h00;
RAM[16'h322D] = 8'h00;
RAM[16'h322E] = 8'h00;
RAM[16'h322F] = 8'h00;
RAM[16'h3230] = 8'h00;
RAM[16'h3231] = 8'h00;
RAM[16'h3232] = 8'h00;
RAM[16'h3233] = 8'h00;
RAM[16'h3234] = 8'h00;
RAM[16'h3235] = 8'h00;
RAM[16'h3236] = 8'h00;
RAM[16'h3237] = 8'h00;
RAM[16'h3238] = 8'h00;
RAM[16'h3239] = 8'h00;
RAM[16'h323A] = 8'h00;
RAM[16'h323B] = 8'h00;
RAM[16'h323C] = 8'h00;
RAM[16'h323D] = 8'h00;
RAM[16'h323E] = 8'h00;
RAM[16'h323F] = 8'h00;
RAM[16'h3240] = 8'h00;
RAM[16'h3241] = 8'h00;
RAM[16'h3242] = 8'h00;
RAM[16'h3243] = 8'h00;
RAM[16'h3244] = 8'h00;
RAM[16'h3245] = 8'h00;
RAM[16'h3246] = 8'h00;
RAM[16'h3247] = 8'h00;
RAM[16'h3248] = 8'h00;
RAM[16'h3249] = 8'h00;
RAM[16'h324A] = 8'h00;
RAM[16'h324B] = 8'h00;
RAM[16'h324C] = 8'h00;
RAM[16'h324D] = 8'h00;
RAM[16'h324E] = 8'h00;
RAM[16'h324F] = 8'h00;
RAM[16'h3250] = 8'h00;
RAM[16'h3251] = 8'h00;
RAM[16'h3252] = 8'h00;
RAM[16'h3253] = 8'h00;
RAM[16'h3254] = 8'h00;
RAM[16'h3255] = 8'h00;
RAM[16'h3256] = 8'h00;
RAM[16'h3257] = 8'h00;
RAM[16'h3258] = 8'h00;
RAM[16'h3259] = 8'h00;
RAM[16'h325A] = 8'h00;
RAM[16'h325B] = 8'h00;
RAM[16'h325C] = 8'h00;
RAM[16'h325D] = 8'h00;
RAM[16'h325E] = 8'h00;
RAM[16'h325F] = 8'h00;
RAM[16'h3260] = 8'h00;
RAM[16'h3261] = 8'h00;
RAM[16'h3262] = 8'h00;
RAM[16'h3263] = 8'h00;
RAM[16'h3264] = 8'h00;
RAM[16'h3265] = 8'h00;
RAM[16'h3266] = 8'h00;
RAM[16'h3267] = 8'h00;
RAM[16'h3268] = 8'h00;
RAM[16'h3269] = 8'h00;
RAM[16'h326A] = 8'h00;
RAM[16'h326B] = 8'h00;
RAM[16'h326C] = 8'h00;
RAM[16'h326D] = 8'h00;
RAM[16'h326E] = 8'h00;
RAM[16'h326F] = 8'h00;
RAM[16'h3270] = 8'h00;
RAM[16'h3271] = 8'h00;
RAM[16'h3272] = 8'h00;
RAM[16'h3273] = 8'h00;
RAM[16'h3274] = 8'h00;
RAM[16'h3275] = 8'h00;
RAM[16'h3276] = 8'h00;
RAM[16'h3277] = 8'h00;
RAM[16'h3278] = 8'h00;
RAM[16'h3279] = 8'h00;
RAM[16'h327A] = 8'h00;
RAM[16'h327B] = 8'h00;
RAM[16'h327C] = 8'h00;
RAM[16'h327D] = 8'h00;
RAM[16'h327E] = 8'h00;
RAM[16'h327F] = 8'h00;
RAM[16'h3280] = 8'h00;
RAM[16'h3281] = 8'h00;
RAM[16'h3282] = 8'h00;
RAM[16'h3283] = 8'h00;
RAM[16'h3284] = 8'h00;
RAM[16'h3285] = 8'h00;
RAM[16'h3286] = 8'h00;
RAM[16'h3287] = 8'h00;
RAM[16'h3288] = 8'h00;
RAM[16'h3289] = 8'h00;
RAM[16'h328A] = 8'h00;
RAM[16'h328B] = 8'h00;
RAM[16'h328C] = 8'h00;
RAM[16'h328D] = 8'h00;
RAM[16'h328E] = 8'h00;
RAM[16'h328F] = 8'h00;
RAM[16'h3290] = 8'h00;
RAM[16'h3291] = 8'h00;
RAM[16'h3292] = 8'h00;
RAM[16'h3293] = 8'h00;
RAM[16'h3294] = 8'h00;
RAM[16'h3295] = 8'h00;
RAM[16'h3296] = 8'h00;
RAM[16'h3297] = 8'h00;
RAM[16'h3298] = 8'h00;
RAM[16'h3299] = 8'h00;
RAM[16'h329A] = 8'h00;
RAM[16'h329B] = 8'h00;
RAM[16'h329C] = 8'h00;
RAM[16'h329D] = 8'h00;
RAM[16'h329E] = 8'h00;
RAM[16'h329F] = 8'h00;
RAM[16'h32A0] = 8'h00;
RAM[16'h32A1] = 8'h00;
RAM[16'h32A2] = 8'h00;
RAM[16'h32A3] = 8'h00;
RAM[16'h32A4] = 8'h00;
RAM[16'h32A5] = 8'h00;
RAM[16'h32A6] = 8'h00;
RAM[16'h32A7] = 8'h00;
RAM[16'h32A8] = 8'h00;
RAM[16'h32A9] = 8'h00;
RAM[16'h32AA] = 8'h00;
RAM[16'h32AB] = 8'h00;
RAM[16'h32AC] = 8'h00;
RAM[16'h32AD] = 8'h00;
RAM[16'h32AE] = 8'h00;
RAM[16'h32AF] = 8'h00;
RAM[16'h32B0] = 8'h00;
RAM[16'h32B1] = 8'h00;
RAM[16'h32B2] = 8'h00;
RAM[16'h32B3] = 8'h00;
RAM[16'h32B4] = 8'h00;
RAM[16'h32B5] = 8'h00;
RAM[16'h32B6] = 8'h00;
RAM[16'h32B7] = 8'h00;
RAM[16'h32B8] = 8'h00;
RAM[16'h32B9] = 8'h00;
RAM[16'h32BA] = 8'h00;
RAM[16'h32BB] = 8'h00;
RAM[16'h32BC] = 8'h00;
RAM[16'h32BD] = 8'h00;
RAM[16'h32BE] = 8'h00;
RAM[16'h32BF] = 8'h00;
RAM[16'h32C0] = 8'h00;
RAM[16'h32C1] = 8'h00;
RAM[16'h32C2] = 8'h00;
RAM[16'h32C3] = 8'h00;
RAM[16'h32C4] = 8'h00;
RAM[16'h32C5] = 8'h00;
RAM[16'h32C6] = 8'h00;
RAM[16'h32C7] = 8'h00;
RAM[16'h32C8] = 8'h00;
RAM[16'h32C9] = 8'h00;
RAM[16'h32CA] = 8'h00;
RAM[16'h32CB] = 8'h00;
RAM[16'h32CC] = 8'h00;
RAM[16'h32CD] = 8'h00;
RAM[16'h32CE] = 8'h00;
RAM[16'h32CF] = 8'h00;
RAM[16'h32D0] = 8'h00;
RAM[16'h32D1] = 8'h00;
RAM[16'h32D2] = 8'h00;
RAM[16'h32D3] = 8'h00;
RAM[16'h32D4] = 8'h00;
RAM[16'h32D5] = 8'h00;
RAM[16'h32D6] = 8'h00;
RAM[16'h32D7] = 8'h00;
RAM[16'h32D8] = 8'h00;
RAM[16'h32D9] = 8'h00;
RAM[16'h32DA] = 8'h00;
RAM[16'h32DB] = 8'h00;
RAM[16'h32DC] = 8'h00;
RAM[16'h32DD] = 8'h00;
RAM[16'h32DE] = 8'h00;
RAM[16'h32DF] = 8'h00;
RAM[16'h32E0] = 8'h00;
RAM[16'h32E1] = 8'h00;
RAM[16'h32E2] = 8'h00;
RAM[16'h32E3] = 8'h00;
RAM[16'h32E4] = 8'h00;
RAM[16'h32E5] = 8'h00;
RAM[16'h32E6] = 8'h00;
RAM[16'h32E7] = 8'h00;
RAM[16'h32E8] = 8'h00;
RAM[16'h32E9] = 8'h00;
RAM[16'h32EA] = 8'h00;
RAM[16'h32EB] = 8'h00;
RAM[16'h32EC] = 8'h00;
RAM[16'h32ED] = 8'h00;
RAM[16'h32EE] = 8'h00;
RAM[16'h32EF] = 8'h00;
RAM[16'h32F0] = 8'h00;
RAM[16'h32F1] = 8'h00;
RAM[16'h32F2] = 8'h00;
RAM[16'h32F3] = 8'h00;
RAM[16'h32F4] = 8'h00;
RAM[16'h32F5] = 8'h00;
RAM[16'h32F6] = 8'h00;
RAM[16'h32F7] = 8'h00;
RAM[16'h32F8] = 8'h00;
RAM[16'h32F9] = 8'h00;
RAM[16'h32FA] = 8'h00;
RAM[16'h32FB] = 8'h00;
RAM[16'h32FC] = 8'h00;
RAM[16'h32FD] = 8'h00;
RAM[16'h32FE] = 8'h00;
RAM[16'h32FF] = 8'h00;
RAM[16'h3300] = 8'h00;
RAM[16'h3301] = 8'h00;
RAM[16'h3302] = 8'h00;
RAM[16'h3303] = 8'h00;
RAM[16'h3304] = 8'h00;
RAM[16'h3305] = 8'h00;
RAM[16'h3306] = 8'h00;
RAM[16'h3307] = 8'h00;
RAM[16'h3308] = 8'h00;
RAM[16'h3309] = 8'h00;
RAM[16'h330A] = 8'h00;
RAM[16'h330B] = 8'h00;
RAM[16'h330C] = 8'h00;
RAM[16'h330D] = 8'h00;
RAM[16'h330E] = 8'h00;
RAM[16'h330F] = 8'h00;
RAM[16'h3310] = 8'h00;
RAM[16'h3311] = 8'h00;
RAM[16'h3312] = 8'h00;
RAM[16'h3313] = 8'h00;
RAM[16'h3314] = 8'h00;
RAM[16'h3315] = 8'h00;
RAM[16'h3316] = 8'h00;
RAM[16'h3317] = 8'h00;
RAM[16'h3318] = 8'h00;
RAM[16'h3319] = 8'h00;
RAM[16'h331A] = 8'h00;
RAM[16'h331B] = 8'h00;
RAM[16'h331C] = 8'h00;
RAM[16'h331D] = 8'h00;
RAM[16'h331E] = 8'h00;
RAM[16'h331F] = 8'h00;
RAM[16'h3320] = 8'h00;
RAM[16'h3321] = 8'h00;
RAM[16'h3322] = 8'h00;
RAM[16'h3323] = 8'h00;
RAM[16'h3324] = 8'h00;
RAM[16'h3325] = 8'h00;
RAM[16'h3326] = 8'h00;
RAM[16'h3327] = 8'h00;
RAM[16'h3328] = 8'h00;
RAM[16'h3329] = 8'h00;
RAM[16'h332A] = 8'h00;
RAM[16'h332B] = 8'h00;
RAM[16'h332C] = 8'h00;
RAM[16'h332D] = 8'h00;
RAM[16'h332E] = 8'h00;
RAM[16'h332F] = 8'h00;
RAM[16'h3330] = 8'h00;
RAM[16'h3331] = 8'h00;
RAM[16'h3332] = 8'h00;
RAM[16'h3333] = 8'h00;
RAM[16'h3334] = 8'h00;
RAM[16'h3335] = 8'h00;
RAM[16'h3336] = 8'h00;
RAM[16'h3337] = 8'h00;
RAM[16'h3338] = 8'h00;
RAM[16'h3339] = 8'h00;
RAM[16'h333A] = 8'h00;
RAM[16'h333B] = 8'h00;
RAM[16'h333C] = 8'h00;
RAM[16'h333D] = 8'h00;
RAM[16'h333E] = 8'h00;
RAM[16'h333F] = 8'h00;
RAM[16'h3340] = 8'h00;
RAM[16'h3341] = 8'h00;
RAM[16'h3342] = 8'h00;
RAM[16'h3343] = 8'h00;
RAM[16'h3344] = 8'h00;
RAM[16'h3345] = 8'h00;
RAM[16'h3346] = 8'h00;
RAM[16'h3347] = 8'h00;
RAM[16'h3348] = 8'h00;
RAM[16'h3349] = 8'h00;
RAM[16'h334A] = 8'h00;
RAM[16'h334B] = 8'h00;
RAM[16'h334C] = 8'h00;
RAM[16'h334D] = 8'h00;
RAM[16'h334E] = 8'h00;
RAM[16'h334F] = 8'h00;
RAM[16'h3350] = 8'h00;
RAM[16'h3351] = 8'h00;
RAM[16'h3352] = 8'h00;
RAM[16'h3353] = 8'h00;
RAM[16'h3354] = 8'h00;
RAM[16'h3355] = 8'h00;
RAM[16'h3356] = 8'h00;
RAM[16'h3357] = 8'h00;
RAM[16'h3358] = 8'h00;
RAM[16'h3359] = 8'h00;
RAM[16'h335A] = 8'h00;
RAM[16'h335B] = 8'h00;
RAM[16'h335C] = 8'h00;
RAM[16'h335D] = 8'h00;
RAM[16'h335E] = 8'h00;
RAM[16'h335F] = 8'h00;
RAM[16'h3360] = 8'h00;
RAM[16'h3361] = 8'h00;
RAM[16'h3362] = 8'h00;
RAM[16'h3363] = 8'h00;
RAM[16'h3364] = 8'h00;
RAM[16'h3365] = 8'h00;
RAM[16'h3366] = 8'h00;
RAM[16'h3367] = 8'h00;
RAM[16'h3368] = 8'h00;
RAM[16'h3369] = 8'h00;
RAM[16'h336A] = 8'h00;
RAM[16'h336B] = 8'h00;
RAM[16'h336C] = 8'h00;
RAM[16'h336D] = 8'h00;
RAM[16'h336E] = 8'h00;
RAM[16'h336F] = 8'h00;
RAM[16'h3370] = 8'h00;
RAM[16'h3371] = 8'h00;
RAM[16'h3372] = 8'h00;
RAM[16'h3373] = 8'h00;
RAM[16'h3374] = 8'h00;
RAM[16'h3375] = 8'h00;
RAM[16'h3376] = 8'h00;
RAM[16'h3377] = 8'h00;
RAM[16'h3378] = 8'h00;
RAM[16'h3379] = 8'h00;
RAM[16'h337A] = 8'h00;
RAM[16'h337B] = 8'h00;
RAM[16'h337C] = 8'h00;
RAM[16'h337D] = 8'h00;
RAM[16'h337E] = 8'h00;
RAM[16'h337F] = 8'h00;
RAM[16'h3380] = 8'h00;
RAM[16'h3381] = 8'h00;
RAM[16'h3382] = 8'h00;
RAM[16'h3383] = 8'h00;
RAM[16'h3384] = 8'h00;
RAM[16'h3385] = 8'h00;
RAM[16'h3386] = 8'h00;
RAM[16'h3387] = 8'h00;
RAM[16'h3388] = 8'h00;
RAM[16'h3389] = 8'h00;
RAM[16'h338A] = 8'h00;
RAM[16'h338B] = 8'h00;
RAM[16'h338C] = 8'h00;
RAM[16'h338D] = 8'h00;
RAM[16'h338E] = 8'h00;
RAM[16'h338F] = 8'h00;
RAM[16'h3390] = 8'h00;
RAM[16'h3391] = 8'h00;
RAM[16'h3392] = 8'h00;
RAM[16'h3393] = 8'h00;
RAM[16'h3394] = 8'h00;
RAM[16'h3395] = 8'h00;
RAM[16'h3396] = 8'h00;
RAM[16'h3397] = 8'h00;
RAM[16'h3398] = 8'h00;
RAM[16'h3399] = 8'h00;
RAM[16'h339A] = 8'h00;
RAM[16'h339B] = 8'h00;
RAM[16'h339C] = 8'h00;
RAM[16'h339D] = 8'h00;
RAM[16'h339E] = 8'h00;
RAM[16'h339F] = 8'h00;
RAM[16'h33A0] = 8'h00;
RAM[16'h33A1] = 8'h00;
RAM[16'h33A2] = 8'h00;
RAM[16'h33A3] = 8'h00;
RAM[16'h33A4] = 8'h00;
RAM[16'h33A5] = 8'h00;
RAM[16'h33A6] = 8'h00;
RAM[16'h33A7] = 8'h00;
RAM[16'h33A8] = 8'h00;
RAM[16'h33A9] = 8'h00;
RAM[16'h33AA] = 8'h00;
RAM[16'h33AB] = 8'h00;
RAM[16'h33AC] = 8'h00;
RAM[16'h33AD] = 8'h00;
RAM[16'h33AE] = 8'h00;
RAM[16'h33AF] = 8'h00;
RAM[16'h33B0] = 8'h00;
RAM[16'h33B1] = 8'h00;
RAM[16'h33B2] = 8'h00;
RAM[16'h33B3] = 8'h00;
RAM[16'h33B4] = 8'h00;
RAM[16'h33B5] = 8'h00;
RAM[16'h33B6] = 8'h00;
RAM[16'h33B7] = 8'h00;
RAM[16'h33B8] = 8'h00;
RAM[16'h33B9] = 8'h00;
RAM[16'h33BA] = 8'h00;
RAM[16'h33BB] = 8'h00;
RAM[16'h33BC] = 8'h00;
RAM[16'h33BD] = 8'h00;
RAM[16'h33BE] = 8'h00;
RAM[16'h33BF] = 8'h00;
RAM[16'h33C0] = 8'h00;
RAM[16'h33C1] = 8'h00;
RAM[16'h33C2] = 8'h00;
RAM[16'h33C3] = 8'h00;
RAM[16'h33C4] = 8'h00;
RAM[16'h33C5] = 8'h00;
RAM[16'h33C6] = 8'h00;
RAM[16'h33C7] = 8'h00;
RAM[16'h33C8] = 8'h00;
RAM[16'h33C9] = 8'h00;
RAM[16'h33CA] = 8'h00;
RAM[16'h33CB] = 8'h00;
RAM[16'h33CC] = 8'h00;
RAM[16'h33CD] = 8'h00;
RAM[16'h33CE] = 8'h00;
RAM[16'h33CF] = 8'h00;
RAM[16'h33D0] = 8'h00;
RAM[16'h33D1] = 8'h00;
RAM[16'h33D2] = 8'h00;
RAM[16'h33D3] = 8'h00;
RAM[16'h33D4] = 8'h00;
RAM[16'h33D5] = 8'h00;
RAM[16'h33D6] = 8'h00;
RAM[16'h33D7] = 8'h00;
RAM[16'h33D8] = 8'h00;
RAM[16'h33D9] = 8'h00;
RAM[16'h33DA] = 8'h00;
RAM[16'h33DB] = 8'h00;
RAM[16'h33DC] = 8'h00;
RAM[16'h33DD] = 8'h00;
RAM[16'h33DE] = 8'h00;
RAM[16'h33DF] = 8'h00;
RAM[16'h33E0] = 8'h00;
RAM[16'h33E1] = 8'h00;
RAM[16'h33E2] = 8'h00;
RAM[16'h33E3] = 8'h00;
RAM[16'h33E4] = 8'h00;
RAM[16'h33E5] = 8'h00;
RAM[16'h33E6] = 8'h00;
RAM[16'h33E7] = 8'h00;
RAM[16'h33E8] = 8'h00;
RAM[16'h33E9] = 8'h00;
RAM[16'h33EA] = 8'h00;
RAM[16'h33EB] = 8'h00;
RAM[16'h33EC] = 8'h00;
RAM[16'h33ED] = 8'h00;
RAM[16'h33EE] = 8'h00;
RAM[16'h33EF] = 8'h00;
RAM[16'h33F0] = 8'h00;
RAM[16'h33F1] = 8'h00;
RAM[16'h33F2] = 8'h00;
RAM[16'h33F3] = 8'h00;
RAM[16'h33F4] = 8'h00;
RAM[16'h33F5] = 8'h00;
RAM[16'h33F6] = 8'h00;
RAM[16'h33F7] = 8'h00;
RAM[16'h33F8] = 8'h00;
RAM[16'h33F9] = 8'h00;
RAM[16'h33FA] = 8'h00;
RAM[16'h33FB] = 8'h00;
RAM[16'h33FC] = 8'h00;
RAM[16'h33FD] = 8'h00;
RAM[16'h33FE] = 8'h00;
RAM[16'h33FF] = 8'h00;
RAM[16'h3400] = 8'h00;
RAM[16'h3401] = 8'h00;
RAM[16'h3402] = 8'h00;
RAM[16'h3403] = 8'h00;
RAM[16'h3404] = 8'h00;
RAM[16'h3405] = 8'h00;
RAM[16'h3406] = 8'h00;
RAM[16'h3407] = 8'h00;
RAM[16'h3408] = 8'h00;
RAM[16'h3409] = 8'h00;
RAM[16'h340A] = 8'h00;
RAM[16'h340B] = 8'h00;
RAM[16'h340C] = 8'h00;
RAM[16'h340D] = 8'h00;
RAM[16'h340E] = 8'h00;
RAM[16'h340F] = 8'h00;
RAM[16'h3410] = 8'h00;
RAM[16'h3411] = 8'h00;
RAM[16'h3412] = 8'h00;
RAM[16'h3413] = 8'h00;
RAM[16'h3414] = 8'h00;
RAM[16'h3415] = 8'h00;
RAM[16'h3416] = 8'h00;
RAM[16'h3417] = 8'h00;
RAM[16'h3418] = 8'h00;
RAM[16'h3419] = 8'h00;
RAM[16'h341A] = 8'h00;
RAM[16'h341B] = 8'h00;
RAM[16'h341C] = 8'h00;
RAM[16'h341D] = 8'h00;
RAM[16'h341E] = 8'h00;
RAM[16'h341F] = 8'h00;
RAM[16'h3420] = 8'h00;
RAM[16'h3421] = 8'h00;
RAM[16'h3422] = 8'h00;
RAM[16'h3423] = 8'h00;
RAM[16'h3424] = 8'h00;
RAM[16'h3425] = 8'h00;
RAM[16'h3426] = 8'h00;
RAM[16'h3427] = 8'h00;
RAM[16'h3428] = 8'h00;
RAM[16'h3429] = 8'h00;
RAM[16'h342A] = 8'h00;
RAM[16'h342B] = 8'h00;
RAM[16'h342C] = 8'h00;
RAM[16'h342D] = 8'h00;
RAM[16'h342E] = 8'h00;
RAM[16'h342F] = 8'h00;
RAM[16'h3430] = 8'h00;
RAM[16'h3431] = 8'h00;
RAM[16'h3432] = 8'h00;
RAM[16'h3433] = 8'h00;
RAM[16'h3434] = 8'h00;
RAM[16'h3435] = 8'h00;
RAM[16'h3436] = 8'h00;
RAM[16'h3437] = 8'h00;
RAM[16'h3438] = 8'h00;
RAM[16'h3439] = 8'h00;
RAM[16'h343A] = 8'h00;
RAM[16'h343B] = 8'h00;
RAM[16'h343C] = 8'h00;
RAM[16'h343D] = 8'h00;
RAM[16'h343E] = 8'h00;
RAM[16'h343F] = 8'h00;
RAM[16'h3440] = 8'h00;
RAM[16'h3441] = 8'h00;
RAM[16'h3442] = 8'h00;
RAM[16'h3443] = 8'h00;
RAM[16'h3444] = 8'h00;
RAM[16'h3445] = 8'h00;
RAM[16'h3446] = 8'h00;
RAM[16'h3447] = 8'h00;
RAM[16'h3448] = 8'h00;
RAM[16'h3449] = 8'h00;
RAM[16'h344A] = 8'h00;
RAM[16'h344B] = 8'h00;
RAM[16'h344C] = 8'h00;
RAM[16'h344D] = 8'h00;
RAM[16'h344E] = 8'h00;
RAM[16'h344F] = 8'h00;
RAM[16'h3450] = 8'h00;
RAM[16'h3451] = 8'h00;
RAM[16'h3452] = 8'h00;
RAM[16'h3453] = 8'h00;
RAM[16'h3454] = 8'h00;
RAM[16'h3455] = 8'h00;
RAM[16'h3456] = 8'h00;
RAM[16'h3457] = 8'h00;
RAM[16'h3458] = 8'h00;
RAM[16'h3459] = 8'h00;
RAM[16'h345A] = 8'h00;
RAM[16'h345B] = 8'h00;
RAM[16'h345C] = 8'h00;
RAM[16'h345D] = 8'h00;
RAM[16'h345E] = 8'h00;
RAM[16'h345F] = 8'h00;
RAM[16'h3460] = 8'h00;
RAM[16'h3461] = 8'h00;
RAM[16'h3462] = 8'h00;
RAM[16'h3463] = 8'h00;
RAM[16'h3464] = 8'h00;
RAM[16'h3465] = 8'h00;
RAM[16'h3466] = 8'h00;
RAM[16'h3467] = 8'h00;
RAM[16'h3468] = 8'h00;
RAM[16'h3469] = 8'h00;
RAM[16'h346A] = 8'h00;
RAM[16'h346B] = 8'h00;
RAM[16'h346C] = 8'h00;
RAM[16'h346D] = 8'h00;
RAM[16'h346E] = 8'h00;
RAM[16'h346F] = 8'h00;
RAM[16'h3470] = 8'h00;
RAM[16'h3471] = 8'h00;
RAM[16'h3472] = 8'h00;
RAM[16'h3473] = 8'h00;
RAM[16'h3474] = 8'h00;
RAM[16'h3475] = 8'h00;
RAM[16'h3476] = 8'h00;
RAM[16'h3477] = 8'h00;
RAM[16'h3478] = 8'h00;
RAM[16'h3479] = 8'h00;
RAM[16'h347A] = 8'h00;
RAM[16'h347B] = 8'h00;
RAM[16'h347C] = 8'h00;
RAM[16'h347D] = 8'h00;
RAM[16'h347E] = 8'h00;
RAM[16'h347F] = 8'h00;
RAM[16'h3480] = 8'h00;
RAM[16'h3481] = 8'h00;
RAM[16'h3482] = 8'h00;
RAM[16'h3483] = 8'h00;
RAM[16'h3484] = 8'h00;
RAM[16'h3485] = 8'h00;
RAM[16'h3486] = 8'h00;
RAM[16'h3487] = 8'h00;
RAM[16'h3488] = 8'h00;
RAM[16'h3489] = 8'h00;
RAM[16'h348A] = 8'h00;
RAM[16'h348B] = 8'h00;
RAM[16'h348C] = 8'h00;
RAM[16'h348D] = 8'h00;
RAM[16'h348E] = 8'h00;
RAM[16'h348F] = 8'h00;
RAM[16'h3490] = 8'h00;
RAM[16'h3491] = 8'h00;
RAM[16'h3492] = 8'h00;
RAM[16'h3493] = 8'h00;
RAM[16'h3494] = 8'h00;
RAM[16'h3495] = 8'h00;
RAM[16'h3496] = 8'h00;
RAM[16'h3497] = 8'h00;
RAM[16'h3498] = 8'h00;
RAM[16'h3499] = 8'h00;
RAM[16'h349A] = 8'h00;
RAM[16'h349B] = 8'h00;
RAM[16'h349C] = 8'h00;
RAM[16'h349D] = 8'h00;
RAM[16'h349E] = 8'h00;
RAM[16'h349F] = 8'h00;
RAM[16'h34A0] = 8'h00;
RAM[16'h34A1] = 8'h00;
RAM[16'h34A2] = 8'h00;
RAM[16'h34A3] = 8'h00;
RAM[16'h34A4] = 8'h00;
RAM[16'h34A5] = 8'h00;
RAM[16'h34A6] = 8'h00;
RAM[16'h34A7] = 8'h00;
RAM[16'h34A8] = 8'h00;
RAM[16'h34A9] = 8'h00;
RAM[16'h34AA] = 8'h00;
RAM[16'h34AB] = 8'h00;
RAM[16'h34AC] = 8'h00;
RAM[16'h34AD] = 8'h00;
RAM[16'h34AE] = 8'h00;
RAM[16'h34AF] = 8'h00;
RAM[16'h34B0] = 8'h00;
RAM[16'h34B1] = 8'h00;
RAM[16'h34B2] = 8'h00;
RAM[16'h34B3] = 8'h00;
RAM[16'h34B4] = 8'h00;
RAM[16'h34B5] = 8'h00;
RAM[16'h34B6] = 8'h00;
RAM[16'h34B7] = 8'h00;
RAM[16'h34B8] = 8'h00;
RAM[16'h34B9] = 8'h00;
RAM[16'h34BA] = 8'h00;
RAM[16'h34BB] = 8'h00;
RAM[16'h34BC] = 8'h00;
RAM[16'h34BD] = 8'h00;
RAM[16'h34BE] = 8'h00;
RAM[16'h34BF] = 8'h00;
RAM[16'h34C0] = 8'h00;
RAM[16'h34C1] = 8'h00;
RAM[16'h34C2] = 8'h00;
RAM[16'h34C3] = 8'h00;
RAM[16'h34C4] = 8'h00;
RAM[16'h34C5] = 8'h00;
RAM[16'h34C6] = 8'h00;
RAM[16'h34C7] = 8'h00;
RAM[16'h34C8] = 8'h00;
RAM[16'h34C9] = 8'h00;
RAM[16'h34CA] = 8'h00;
RAM[16'h34CB] = 8'h00;
RAM[16'h34CC] = 8'h00;
RAM[16'h34CD] = 8'h00;
RAM[16'h34CE] = 8'h00;
RAM[16'h34CF] = 8'h00;
RAM[16'h34D0] = 8'h00;
RAM[16'h34D1] = 8'h00;
RAM[16'h34D2] = 8'h00;
RAM[16'h34D3] = 8'h00;
RAM[16'h34D4] = 8'h00;
RAM[16'h34D5] = 8'h00;
RAM[16'h34D6] = 8'h00;
RAM[16'h34D7] = 8'h00;
RAM[16'h34D8] = 8'h00;
RAM[16'h34D9] = 8'h00;
RAM[16'h34DA] = 8'h00;
RAM[16'h34DB] = 8'h00;
RAM[16'h34DC] = 8'h00;
RAM[16'h34DD] = 8'h00;
RAM[16'h34DE] = 8'h00;
RAM[16'h34DF] = 8'h00;
RAM[16'h34E0] = 8'h00;
RAM[16'h34E1] = 8'h00;
RAM[16'h34E2] = 8'h00;
RAM[16'h34E3] = 8'h00;
RAM[16'h34E4] = 8'h00;
RAM[16'h34E5] = 8'h00;
RAM[16'h34E6] = 8'h00;
RAM[16'h34E7] = 8'h00;
RAM[16'h34E8] = 8'h00;
RAM[16'h34E9] = 8'h00;
RAM[16'h34EA] = 8'h00;
RAM[16'h34EB] = 8'h00;
RAM[16'h34EC] = 8'h00;
RAM[16'h34ED] = 8'h00;
RAM[16'h34EE] = 8'h00;
RAM[16'h34EF] = 8'h00;
RAM[16'h34F0] = 8'h00;
RAM[16'h34F1] = 8'h00;
RAM[16'h34F2] = 8'h00;
RAM[16'h34F3] = 8'h00;
RAM[16'h34F4] = 8'h00;
RAM[16'h34F5] = 8'h00;
RAM[16'h34F6] = 8'h00;
RAM[16'h34F7] = 8'h00;
RAM[16'h34F8] = 8'h00;
RAM[16'h34F9] = 8'h00;
RAM[16'h34FA] = 8'h00;
RAM[16'h34FB] = 8'h00;
RAM[16'h34FC] = 8'h00;
RAM[16'h34FD] = 8'h00;
RAM[16'h34FE] = 8'h00;
RAM[16'h34FF] = 8'h00;
RAM[16'h3500] = 8'h00;
RAM[16'h3501] = 8'h00;
RAM[16'h3502] = 8'h00;
RAM[16'h3503] = 8'h00;
RAM[16'h3504] = 8'h00;
RAM[16'h3505] = 8'h00;
RAM[16'h3506] = 8'h00;
RAM[16'h3507] = 8'h00;
RAM[16'h3508] = 8'h00;
RAM[16'h3509] = 8'h00;
RAM[16'h350A] = 8'h00;
RAM[16'h350B] = 8'h00;
RAM[16'h350C] = 8'h00;
RAM[16'h350D] = 8'h00;
RAM[16'h350E] = 8'h00;
RAM[16'h350F] = 8'h00;
RAM[16'h3510] = 8'h00;
RAM[16'h3511] = 8'h00;
RAM[16'h3512] = 8'h00;
RAM[16'h3513] = 8'h00;
RAM[16'h3514] = 8'h00;
RAM[16'h3515] = 8'h00;
RAM[16'h3516] = 8'h00;
RAM[16'h3517] = 8'h00;
RAM[16'h3518] = 8'h00;
RAM[16'h3519] = 8'h00;
RAM[16'h351A] = 8'h00;
RAM[16'h351B] = 8'h00;
RAM[16'h351C] = 8'h00;
RAM[16'h351D] = 8'h00;
RAM[16'h351E] = 8'h00;
RAM[16'h351F] = 8'h00;
RAM[16'h3520] = 8'h00;
RAM[16'h3521] = 8'h00;
RAM[16'h3522] = 8'h00;
RAM[16'h3523] = 8'h00;
RAM[16'h3524] = 8'h00;
RAM[16'h3525] = 8'h00;
RAM[16'h3526] = 8'h00;
RAM[16'h3527] = 8'h00;
RAM[16'h3528] = 8'h00;
RAM[16'h3529] = 8'h00;
RAM[16'h352A] = 8'h00;
RAM[16'h352B] = 8'h00;
RAM[16'h352C] = 8'h00;
RAM[16'h352D] = 8'h00;
RAM[16'h352E] = 8'h00;
RAM[16'h352F] = 8'h00;
RAM[16'h3530] = 8'h00;
RAM[16'h3531] = 8'h00;
RAM[16'h3532] = 8'h00;
RAM[16'h3533] = 8'h00;
RAM[16'h3534] = 8'h00;
RAM[16'h3535] = 8'h00;
RAM[16'h3536] = 8'h00;
RAM[16'h3537] = 8'h00;
RAM[16'h3538] = 8'h00;
RAM[16'h3539] = 8'h00;
RAM[16'h353A] = 8'h00;
RAM[16'h353B] = 8'h00;
RAM[16'h353C] = 8'h00;
RAM[16'h353D] = 8'h00;
RAM[16'h353E] = 8'h00;
RAM[16'h353F] = 8'h00;
RAM[16'h3540] = 8'h00;
RAM[16'h3541] = 8'h00;
RAM[16'h3542] = 8'h00;
RAM[16'h3543] = 8'h00;
RAM[16'h3544] = 8'h00;
RAM[16'h3545] = 8'h00;
RAM[16'h3546] = 8'h00;
RAM[16'h3547] = 8'h00;
RAM[16'h3548] = 8'h00;
RAM[16'h3549] = 8'h00;
RAM[16'h354A] = 8'h00;
RAM[16'h354B] = 8'h00;
RAM[16'h354C] = 8'h00;
RAM[16'h354D] = 8'h00;
RAM[16'h354E] = 8'h00;
RAM[16'h354F] = 8'h00;
RAM[16'h3550] = 8'h00;
RAM[16'h3551] = 8'h00;
RAM[16'h3552] = 8'h00;
RAM[16'h3553] = 8'h00;
RAM[16'h3554] = 8'h00;
RAM[16'h3555] = 8'h00;
RAM[16'h3556] = 8'h00;
RAM[16'h3557] = 8'h00;
RAM[16'h3558] = 8'h00;
RAM[16'h3559] = 8'h00;
RAM[16'h355A] = 8'h00;
RAM[16'h355B] = 8'h00;
RAM[16'h355C] = 8'h00;
RAM[16'h355D] = 8'h00;
RAM[16'h355E] = 8'h00;
RAM[16'h355F] = 8'h00;
RAM[16'h3560] = 8'h00;
RAM[16'h3561] = 8'h00;
RAM[16'h3562] = 8'h00;
RAM[16'h3563] = 8'h00;
RAM[16'h3564] = 8'h00;
RAM[16'h3565] = 8'h00;
RAM[16'h3566] = 8'h00;
RAM[16'h3567] = 8'h00;
RAM[16'h3568] = 8'h00;
RAM[16'h3569] = 8'h00;
RAM[16'h356A] = 8'h00;
RAM[16'h356B] = 8'h00;
RAM[16'h356C] = 8'h00;
RAM[16'h356D] = 8'h00;
RAM[16'h356E] = 8'h00;
RAM[16'h356F] = 8'h00;
RAM[16'h3570] = 8'h00;
RAM[16'h3571] = 8'h00;
RAM[16'h3572] = 8'h00;
RAM[16'h3573] = 8'h00;
RAM[16'h3574] = 8'h00;
RAM[16'h3575] = 8'h00;
RAM[16'h3576] = 8'h00;
RAM[16'h3577] = 8'h00;
RAM[16'h3578] = 8'h00;
RAM[16'h3579] = 8'h00;
RAM[16'h357A] = 8'h00;
RAM[16'h357B] = 8'h00;
RAM[16'h357C] = 8'h00;
RAM[16'h357D] = 8'h00;
RAM[16'h357E] = 8'h00;
RAM[16'h357F] = 8'h00;
RAM[16'h3580] = 8'h00;
RAM[16'h3581] = 8'h00;
RAM[16'h3582] = 8'h00;
RAM[16'h3583] = 8'h00;
RAM[16'h3584] = 8'h00;
RAM[16'h3585] = 8'h00;
RAM[16'h3586] = 8'h00;
RAM[16'h3587] = 8'h00;
RAM[16'h3588] = 8'h00;
RAM[16'h3589] = 8'h00;
RAM[16'h358A] = 8'h00;
RAM[16'h358B] = 8'h00;
RAM[16'h358C] = 8'h00;
RAM[16'h358D] = 8'h00;
RAM[16'h358E] = 8'h00;
RAM[16'h358F] = 8'h00;
RAM[16'h3590] = 8'h00;
RAM[16'h3591] = 8'h00;
RAM[16'h3592] = 8'h00;
RAM[16'h3593] = 8'h00;
RAM[16'h3594] = 8'h00;
RAM[16'h3595] = 8'h00;
RAM[16'h3596] = 8'h00;
RAM[16'h3597] = 8'h00;
RAM[16'h3598] = 8'h00;
RAM[16'h3599] = 8'h00;
RAM[16'h359A] = 8'h00;
RAM[16'h359B] = 8'h00;
RAM[16'h359C] = 8'h00;
RAM[16'h359D] = 8'h00;
RAM[16'h359E] = 8'h00;
RAM[16'h359F] = 8'h00;
RAM[16'h35A0] = 8'h00;
RAM[16'h35A1] = 8'h00;
RAM[16'h35A2] = 8'h00;
RAM[16'h35A3] = 8'h00;
RAM[16'h35A4] = 8'h00;
RAM[16'h35A5] = 8'h00;
RAM[16'h35A6] = 8'h00;
RAM[16'h35A7] = 8'h00;
RAM[16'h35A8] = 8'h00;
RAM[16'h35A9] = 8'h00;
RAM[16'h35AA] = 8'h00;
RAM[16'h35AB] = 8'h00;
RAM[16'h35AC] = 8'h00;
RAM[16'h35AD] = 8'h00;
RAM[16'h35AE] = 8'h00;
RAM[16'h35AF] = 8'h00;
RAM[16'h35B0] = 8'h00;
RAM[16'h35B1] = 8'h00;
RAM[16'h35B2] = 8'h00;
RAM[16'h35B3] = 8'h00;
RAM[16'h35B4] = 8'h00;
RAM[16'h35B5] = 8'h00;
RAM[16'h35B6] = 8'h00;
RAM[16'h35B7] = 8'h00;
RAM[16'h35B8] = 8'h00;
RAM[16'h35B9] = 8'h00;
RAM[16'h35BA] = 8'h00;
RAM[16'h35BB] = 8'h00;
RAM[16'h35BC] = 8'h00;
RAM[16'h35BD] = 8'h00;
RAM[16'h35BE] = 8'h00;
RAM[16'h35BF] = 8'h00;
RAM[16'h35C0] = 8'h00;
RAM[16'h35C1] = 8'h00;
RAM[16'h35C2] = 8'h00;
RAM[16'h35C3] = 8'h00;
RAM[16'h35C4] = 8'h00;
RAM[16'h35C5] = 8'h00;
RAM[16'h35C6] = 8'h00;
RAM[16'h35C7] = 8'h00;
RAM[16'h35C8] = 8'h00;
RAM[16'h35C9] = 8'h00;
RAM[16'h35CA] = 8'h00;
RAM[16'h35CB] = 8'h00;
RAM[16'h35CC] = 8'h00;
RAM[16'h35CD] = 8'h00;
RAM[16'h35CE] = 8'h00;
RAM[16'h35CF] = 8'h00;
RAM[16'h35D0] = 8'h00;
RAM[16'h35D1] = 8'h00;
RAM[16'h35D2] = 8'h00;
RAM[16'h35D3] = 8'h00;
RAM[16'h35D4] = 8'h00;
RAM[16'h35D5] = 8'h00;
RAM[16'h35D6] = 8'h00;
RAM[16'h35D7] = 8'h00;
RAM[16'h35D8] = 8'h00;
RAM[16'h35D9] = 8'h00;
RAM[16'h35DA] = 8'h00;
RAM[16'h35DB] = 8'h00;
RAM[16'h35DC] = 8'h00;
RAM[16'h35DD] = 8'h00;
RAM[16'h35DE] = 8'h00;
RAM[16'h35DF] = 8'h00;
RAM[16'h35E0] = 8'h00;
RAM[16'h35E1] = 8'h00;
RAM[16'h35E2] = 8'h00;
RAM[16'h35E3] = 8'h00;
RAM[16'h35E4] = 8'h00;
RAM[16'h35E5] = 8'h00;
RAM[16'h35E6] = 8'h00;
RAM[16'h35E7] = 8'h00;
RAM[16'h35E8] = 8'h00;
RAM[16'h35E9] = 8'h00;
RAM[16'h35EA] = 8'h00;
RAM[16'h35EB] = 8'h00;
RAM[16'h35EC] = 8'h00;
RAM[16'h35ED] = 8'h00;
RAM[16'h35EE] = 8'h00;
RAM[16'h35EF] = 8'h00;
RAM[16'h35F0] = 8'h00;
RAM[16'h35F1] = 8'h00;
RAM[16'h35F2] = 8'h00;
RAM[16'h35F3] = 8'h00;
RAM[16'h35F4] = 8'h00;
RAM[16'h35F5] = 8'h00;
RAM[16'h35F6] = 8'h00;
RAM[16'h35F7] = 8'h00;
RAM[16'h35F8] = 8'h00;
RAM[16'h35F9] = 8'h00;
RAM[16'h35FA] = 8'h00;
RAM[16'h35FB] = 8'h00;
RAM[16'h35FC] = 8'h00;
RAM[16'h35FD] = 8'h00;
RAM[16'h35FE] = 8'h00;
RAM[16'h35FF] = 8'h00;
RAM[16'h3600] = 8'h00;
RAM[16'h3601] = 8'h00;
RAM[16'h3602] = 8'h00;
RAM[16'h3603] = 8'h00;
RAM[16'h3604] = 8'h00;
RAM[16'h3605] = 8'h00;
RAM[16'h3606] = 8'h00;
RAM[16'h3607] = 8'h00;
RAM[16'h3608] = 8'h00;
RAM[16'h3609] = 8'h00;
RAM[16'h360A] = 8'h00;
RAM[16'h360B] = 8'h00;
RAM[16'h360C] = 8'h00;
RAM[16'h360D] = 8'h00;
RAM[16'h360E] = 8'h00;
RAM[16'h360F] = 8'h00;
RAM[16'h3610] = 8'h00;
RAM[16'h3611] = 8'h00;
RAM[16'h3612] = 8'h00;
RAM[16'h3613] = 8'h00;
RAM[16'h3614] = 8'h00;
RAM[16'h3615] = 8'h00;
RAM[16'h3616] = 8'h00;
RAM[16'h3617] = 8'h00;
RAM[16'h3618] = 8'h00;
RAM[16'h3619] = 8'h00;
RAM[16'h361A] = 8'h00;
RAM[16'h361B] = 8'h00;
RAM[16'h361C] = 8'h00;
RAM[16'h361D] = 8'h00;
RAM[16'h361E] = 8'h00;
RAM[16'h361F] = 8'h00;
RAM[16'h3620] = 8'h00;
RAM[16'h3621] = 8'h00;
RAM[16'h3622] = 8'h00;
RAM[16'h3623] = 8'h00;
RAM[16'h3624] = 8'h00;
RAM[16'h3625] = 8'h00;
RAM[16'h3626] = 8'h00;
RAM[16'h3627] = 8'h00;
RAM[16'h3628] = 8'h00;
RAM[16'h3629] = 8'h00;
RAM[16'h362A] = 8'h00;
RAM[16'h362B] = 8'h00;
RAM[16'h362C] = 8'h00;
RAM[16'h362D] = 8'h00;
RAM[16'h362E] = 8'h00;
RAM[16'h362F] = 8'h00;
RAM[16'h3630] = 8'h00;
RAM[16'h3631] = 8'h00;
RAM[16'h3632] = 8'h00;
RAM[16'h3633] = 8'h00;
RAM[16'h3634] = 8'h00;
RAM[16'h3635] = 8'h00;
RAM[16'h3636] = 8'h00;
RAM[16'h3637] = 8'h00;
RAM[16'h3638] = 8'h00;
RAM[16'h3639] = 8'h00;
RAM[16'h363A] = 8'h00;
RAM[16'h363B] = 8'h00;
RAM[16'h363C] = 8'h00;
RAM[16'h363D] = 8'h00;
RAM[16'h363E] = 8'h00;
RAM[16'h363F] = 8'h00;
RAM[16'h3640] = 8'h00;
RAM[16'h3641] = 8'h00;
RAM[16'h3642] = 8'h00;
RAM[16'h3643] = 8'h00;
RAM[16'h3644] = 8'h00;
RAM[16'h3645] = 8'h00;
RAM[16'h3646] = 8'h00;
RAM[16'h3647] = 8'h00;
RAM[16'h3648] = 8'h00;
RAM[16'h3649] = 8'h00;
RAM[16'h364A] = 8'h00;
RAM[16'h364B] = 8'h00;
RAM[16'h364C] = 8'h00;
RAM[16'h364D] = 8'h00;
RAM[16'h364E] = 8'h00;
RAM[16'h364F] = 8'h00;
RAM[16'h3650] = 8'h00;
RAM[16'h3651] = 8'h00;
RAM[16'h3652] = 8'h00;
RAM[16'h3653] = 8'h00;
RAM[16'h3654] = 8'h00;
RAM[16'h3655] = 8'h00;
RAM[16'h3656] = 8'h00;
RAM[16'h3657] = 8'h00;
RAM[16'h3658] = 8'h00;
RAM[16'h3659] = 8'h00;
RAM[16'h365A] = 8'h00;
RAM[16'h365B] = 8'h00;
RAM[16'h365C] = 8'h00;
RAM[16'h365D] = 8'h00;
RAM[16'h365E] = 8'h00;
RAM[16'h365F] = 8'h00;
RAM[16'h3660] = 8'h00;
RAM[16'h3661] = 8'h00;
RAM[16'h3662] = 8'h00;
RAM[16'h3663] = 8'h00;
RAM[16'h3664] = 8'h00;
RAM[16'h3665] = 8'h00;
RAM[16'h3666] = 8'h00;
RAM[16'h3667] = 8'h00;
RAM[16'h3668] = 8'h00;
RAM[16'h3669] = 8'h00;
RAM[16'h366A] = 8'h00;
RAM[16'h366B] = 8'h00;
RAM[16'h366C] = 8'h00;
RAM[16'h366D] = 8'h00;
RAM[16'h366E] = 8'h00;
RAM[16'h366F] = 8'h00;
RAM[16'h3670] = 8'h00;
RAM[16'h3671] = 8'h00;
RAM[16'h3672] = 8'h00;
RAM[16'h3673] = 8'h00;
RAM[16'h3674] = 8'h00;
RAM[16'h3675] = 8'h00;
RAM[16'h3676] = 8'h00;
RAM[16'h3677] = 8'h00;
RAM[16'h3678] = 8'h00;
RAM[16'h3679] = 8'h00;
RAM[16'h367A] = 8'h00;
RAM[16'h367B] = 8'h00;
RAM[16'h367C] = 8'h00;
RAM[16'h367D] = 8'h00;
RAM[16'h367E] = 8'h00;
RAM[16'h367F] = 8'h00;
RAM[16'h3680] = 8'h00;
RAM[16'h3681] = 8'h00;
RAM[16'h3682] = 8'h00;
RAM[16'h3683] = 8'h00;
RAM[16'h3684] = 8'h00;
RAM[16'h3685] = 8'h00;
RAM[16'h3686] = 8'h00;
RAM[16'h3687] = 8'h00;
RAM[16'h3688] = 8'h00;
RAM[16'h3689] = 8'h00;
RAM[16'h368A] = 8'h00;
RAM[16'h368B] = 8'h00;
RAM[16'h368C] = 8'h00;
RAM[16'h368D] = 8'h00;
RAM[16'h368E] = 8'h00;
RAM[16'h368F] = 8'h00;
RAM[16'h3690] = 8'h00;
RAM[16'h3691] = 8'h00;
RAM[16'h3692] = 8'h00;
RAM[16'h3693] = 8'h00;
RAM[16'h3694] = 8'h00;
RAM[16'h3695] = 8'h00;
RAM[16'h3696] = 8'h00;
RAM[16'h3697] = 8'h00;
RAM[16'h3698] = 8'h00;
RAM[16'h3699] = 8'h00;
RAM[16'h369A] = 8'h00;
RAM[16'h369B] = 8'h00;
RAM[16'h369C] = 8'h00;
RAM[16'h369D] = 8'h00;
RAM[16'h369E] = 8'h00;
RAM[16'h369F] = 8'h00;
RAM[16'h36A0] = 8'h00;
RAM[16'h36A1] = 8'h00;
RAM[16'h36A2] = 8'h00;
RAM[16'h36A3] = 8'h00;
RAM[16'h36A4] = 8'h00;
RAM[16'h36A5] = 8'h00;
RAM[16'h36A6] = 8'h00;
RAM[16'h36A7] = 8'h00;
RAM[16'h36A8] = 8'h00;
RAM[16'h36A9] = 8'h00;
RAM[16'h36AA] = 8'h00;
RAM[16'h36AB] = 8'h00;
RAM[16'h36AC] = 8'h00;
RAM[16'h36AD] = 8'h00;
RAM[16'h36AE] = 8'h00;
RAM[16'h36AF] = 8'h00;
RAM[16'h36B0] = 8'h00;
RAM[16'h36B1] = 8'h00;
RAM[16'h36B2] = 8'h00;
RAM[16'h36B3] = 8'h00;
RAM[16'h36B4] = 8'h00;
RAM[16'h36B5] = 8'h00;
RAM[16'h36B6] = 8'h00;
RAM[16'h36B7] = 8'h00;
RAM[16'h36B8] = 8'h00;
RAM[16'h36B9] = 8'h00;
RAM[16'h36BA] = 8'h00;
RAM[16'h36BB] = 8'h00;
RAM[16'h36BC] = 8'h00;
RAM[16'h36BD] = 8'h00;
RAM[16'h36BE] = 8'h00;
RAM[16'h36BF] = 8'h00;
RAM[16'h36C0] = 8'h00;
RAM[16'h36C1] = 8'h00;
RAM[16'h36C2] = 8'h00;
RAM[16'h36C3] = 8'h00;
RAM[16'h36C4] = 8'h00;
RAM[16'h36C5] = 8'h00;
RAM[16'h36C6] = 8'h00;
RAM[16'h36C7] = 8'h00;
RAM[16'h36C8] = 8'h00;
RAM[16'h36C9] = 8'h00;
RAM[16'h36CA] = 8'h00;
RAM[16'h36CB] = 8'h00;
RAM[16'h36CC] = 8'h00;
RAM[16'h36CD] = 8'h00;
RAM[16'h36CE] = 8'h00;
RAM[16'h36CF] = 8'h00;
RAM[16'h36D0] = 8'h00;
RAM[16'h36D1] = 8'h00;
RAM[16'h36D2] = 8'h00;
RAM[16'h36D3] = 8'h00;
RAM[16'h36D4] = 8'h00;
RAM[16'h36D5] = 8'h00;
RAM[16'h36D6] = 8'h00;
RAM[16'h36D7] = 8'h00;
RAM[16'h36D8] = 8'h00;
RAM[16'h36D9] = 8'h00;
RAM[16'h36DA] = 8'h00;
RAM[16'h36DB] = 8'h00;
RAM[16'h36DC] = 8'h00;
RAM[16'h36DD] = 8'h00;
RAM[16'h36DE] = 8'h00;
RAM[16'h36DF] = 8'h00;
RAM[16'h36E0] = 8'h00;
RAM[16'h36E1] = 8'h00;
RAM[16'h36E2] = 8'h00;
RAM[16'h36E3] = 8'h00;
RAM[16'h36E4] = 8'h00;
RAM[16'h36E5] = 8'h00;
RAM[16'h36E6] = 8'h00;
RAM[16'h36E7] = 8'h00;
RAM[16'h36E8] = 8'h00;
RAM[16'h36E9] = 8'h00;
RAM[16'h36EA] = 8'h00;
RAM[16'h36EB] = 8'h00;
RAM[16'h36EC] = 8'h00;
RAM[16'h36ED] = 8'h00;
RAM[16'h36EE] = 8'h00;
RAM[16'h36EF] = 8'h00;
RAM[16'h36F0] = 8'h00;
RAM[16'h36F1] = 8'h00;
RAM[16'h36F2] = 8'h00;
RAM[16'h36F3] = 8'h00;
RAM[16'h36F4] = 8'h00;
RAM[16'h36F5] = 8'h00;
RAM[16'h36F6] = 8'h00;
RAM[16'h36F7] = 8'h00;
RAM[16'h36F8] = 8'h00;
RAM[16'h36F9] = 8'h00;
RAM[16'h36FA] = 8'h00;
RAM[16'h36FB] = 8'h00;
RAM[16'h36FC] = 8'h00;
RAM[16'h36FD] = 8'h00;
RAM[16'h36FE] = 8'h00;
RAM[16'h36FF] = 8'h00;
RAM[16'h3700] = 8'h00;
RAM[16'h3701] = 8'h00;
RAM[16'h3702] = 8'h00;
RAM[16'h3703] = 8'h00;
RAM[16'h3704] = 8'h00;
RAM[16'h3705] = 8'h00;
RAM[16'h3706] = 8'h00;
RAM[16'h3707] = 8'h00;
RAM[16'h3708] = 8'h00;
RAM[16'h3709] = 8'h00;
RAM[16'h370A] = 8'h00;
RAM[16'h370B] = 8'h00;
RAM[16'h370C] = 8'h00;
RAM[16'h370D] = 8'h00;
RAM[16'h370E] = 8'h00;
RAM[16'h370F] = 8'h00;
RAM[16'h3710] = 8'h00;
RAM[16'h3711] = 8'h00;
RAM[16'h3712] = 8'h00;
RAM[16'h3713] = 8'h00;
RAM[16'h3714] = 8'h00;
RAM[16'h3715] = 8'h00;
RAM[16'h3716] = 8'h00;
RAM[16'h3717] = 8'h00;
RAM[16'h3718] = 8'h00;
RAM[16'h3719] = 8'h00;
RAM[16'h371A] = 8'h00;
RAM[16'h371B] = 8'h00;
RAM[16'h371C] = 8'h00;
RAM[16'h371D] = 8'h00;
RAM[16'h371E] = 8'h00;
RAM[16'h371F] = 8'h00;
RAM[16'h3720] = 8'h00;
RAM[16'h3721] = 8'h00;
RAM[16'h3722] = 8'h00;
RAM[16'h3723] = 8'h00;
RAM[16'h3724] = 8'h00;
RAM[16'h3725] = 8'h00;
RAM[16'h3726] = 8'h00;
RAM[16'h3727] = 8'h00;
RAM[16'h3728] = 8'h00;
RAM[16'h3729] = 8'h00;
RAM[16'h372A] = 8'h00;
RAM[16'h372B] = 8'h00;
RAM[16'h372C] = 8'h00;
RAM[16'h372D] = 8'h00;
RAM[16'h372E] = 8'h00;
RAM[16'h372F] = 8'h00;
RAM[16'h3730] = 8'h00;
RAM[16'h3731] = 8'h00;
RAM[16'h3732] = 8'h00;
RAM[16'h3733] = 8'h00;
RAM[16'h3734] = 8'h00;
RAM[16'h3735] = 8'h00;
RAM[16'h3736] = 8'h00;
RAM[16'h3737] = 8'h00;
RAM[16'h3738] = 8'h00;
RAM[16'h3739] = 8'h00;
RAM[16'h373A] = 8'h00;
RAM[16'h373B] = 8'h00;
RAM[16'h373C] = 8'h00;
RAM[16'h373D] = 8'h00;
RAM[16'h373E] = 8'h00;
RAM[16'h373F] = 8'h00;
RAM[16'h3740] = 8'h00;
RAM[16'h3741] = 8'h00;
RAM[16'h3742] = 8'h00;
RAM[16'h3743] = 8'h00;
RAM[16'h3744] = 8'h00;
RAM[16'h3745] = 8'h00;
RAM[16'h3746] = 8'h00;
RAM[16'h3747] = 8'h00;
RAM[16'h3748] = 8'h00;
RAM[16'h3749] = 8'h00;
RAM[16'h374A] = 8'h00;
RAM[16'h374B] = 8'h00;
RAM[16'h374C] = 8'h00;
RAM[16'h374D] = 8'h00;
RAM[16'h374E] = 8'h00;
RAM[16'h374F] = 8'h00;
RAM[16'h3750] = 8'h00;
RAM[16'h3751] = 8'h00;
RAM[16'h3752] = 8'h00;
RAM[16'h3753] = 8'h00;
RAM[16'h3754] = 8'h00;
RAM[16'h3755] = 8'h00;
RAM[16'h3756] = 8'h00;
RAM[16'h3757] = 8'h00;
RAM[16'h3758] = 8'h00;
RAM[16'h3759] = 8'h00;
RAM[16'h375A] = 8'h00;
RAM[16'h375B] = 8'h00;
RAM[16'h375C] = 8'h00;
RAM[16'h375D] = 8'h00;
RAM[16'h375E] = 8'h00;
RAM[16'h375F] = 8'h00;
RAM[16'h3760] = 8'h00;
RAM[16'h3761] = 8'h00;
RAM[16'h3762] = 8'h00;
RAM[16'h3763] = 8'h00;
RAM[16'h3764] = 8'h00;
RAM[16'h3765] = 8'h00;
RAM[16'h3766] = 8'h00;
RAM[16'h3767] = 8'h00;
RAM[16'h3768] = 8'h00;
RAM[16'h3769] = 8'h00;
RAM[16'h376A] = 8'h00;
RAM[16'h376B] = 8'h00;
RAM[16'h376C] = 8'h00;
RAM[16'h376D] = 8'h00;
RAM[16'h376E] = 8'h00;
RAM[16'h376F] = 8'h00;
RAM[16'h3770] = 8'h00;
RAM[16'h3771] = 8'h00;
RAM[16'h3772] = 8'h00;
RAM[16'h3773] = 8'h00;
RAM[16'h3774] = 8'h00;
RAM[16'h3775] = 8'h00;
RAM[16'h3776] = 8'h00;
RAM[16'h3777] = 8'h00;
RAM[16'h3778] = 8'h00;
RAM[16'h3779] = 8'h00;
RAM[16'h377A] = 8'h00;
RAM[16'h377B] = 8'h00;
RAM[16'h377C] = 8'h00;
RAM[16'h377D] = 8'h00;
RAM[16'h377E] = 8'h00;
RAM[16'h377F] = 8'h00;
RAM[16'h3780] = 8'h00;
RAM[16'h3781] = 8'h00;
RAM[16'h3782] = 8'h00;
RAM[16'h3783] = 8'h00;
RAM[16'h3784] = 8'h00;
RAM[16'h3785] = 8'h00;
RAM[16'h3786] = 8'h00;
RAM[16'h3787] = 8'h00;
RAM[16'h3788] = 8'h00;
RAM[16'h3789] = 8'h00;
RAM[16'h378A] = 8'h00;
RAM[16'h378B] = 8'h00;
RAM[16'h378C] = 8'h00;
RAM[16'h378D] = 8'h00;
RAM[16'h378E] = 8'h00;
RAM[16'h378F] = 8'h00;
RAM[16'h3790] = 8'h00;
RAM[16'h3791] = 8'h00;
RAM[16'h3792] = 8'h00;
RAM[16'h3793] = 8'h00;
RAM[16'h3794] = 8'h00;
RAM[16'h3795] = 8'h00;
RAM[16'h3796] = 8'h00;
RAM[16'h3797] = 8'h00;
RAM[16'h3798] = 8'h00;
RAM[16'h3799] = 8'h00;
RAM[16'h379A] = 8'h00;
RAM[16'h379B] = 8'h00;
RAM[16'h379C] = 8'h00;
RAM[16'h379D] = 8'h00;
RAM[16'h379E] = 8'h00;
RAM[16'h379F] = 8'h00;
RAM[16'h37A0] = 8'h00;
RAM[16'h37A1] = 8'h00;
RAM[16'h37A2] = 8'h00;
RAM[16'h37A3] = 8'h00;
RAM[16'h37A4] = 8'h00;
RAM[16'h37A5] = 8'h00;
RAM[16'h37A6] = 8'h00;
RAM[16'h37A7] = 8'h00;
RAM[16'h37A8] = 8'h00;
RAM[16'h37A9] = 8'h00;
RAM[16'h37AA] = 8'h00;
RAM[16'h37AB] = 8'h00;
RAM[16'h37AC] = 8'h00;
RAM[16'h37AD] = 8'h00;
RAM[16'h37AE] = 8'h00;
RAM[16'h37AF] = 8'h00;
RAM[16'h37B0] = 8'h00;
RAM[16'h37B1] = 8'h00;
RAM[16'h37B2] = 8'h00;
RAM[16'h37B3] = 8'h00;
RAM[16'h37B4] = 8'h00;
RAM[16'h37B5] = 8'h00;
RAM[16'h37B6] = 8'h00;
RAM[16'h37B7] = 8'h00;
RAM[16'h37B8] = 8'h00;
RAM[16'h37B9] = 8'h00;
RAM[16'h37BA] = 8'h00;
RAM[16'h37BB] = 8'h00;
RAM[16'h37BC] = 8'h00;
RAM[16'h37BD] = 8'h00;
RAM[16'h37BE] = 8'h00;
RAM[16'h37BF] = 8'h00;
RAM[16'h37C0] = 8'h00;
RAM[16'h37C1] = 8'h00;
RAM[16'h37C2] = 8'h00;
RAM[16'h37C3] = 8'h00;
RAM[16'h37C4] = 8'h00;
RAM[16'h37C5] = 8'h00;
RAM[16'h37C6] = 8'h00;
RAM[16'h37C7] = 8'h00;
RAM[16'h37C8] = 8'h00;
RAM[16'h37C9] = 8'h00;
RAM[16'h37CA] = 8'h00;
RAM[16'h37CB] = 8'h00;
RAM[16'h37CC] = 8'h00;
RAM[16'h37CD] = 8'h00;
RAM[16'h37CE] = 8'h00;
RAM[16'h37CF] = 8'h00;
RAM[16'h37D0] = 8'h00;
RAM[16'h37D1] = 8'h00;
RAM[16'h37D2] = 8'h00;
RAM[16'h37D3] = 8'h00;
RAM[16'h37D4] = 8'h00;
RAM[16'h37D5] = 8'h00;
RAM[16'h37D6] = 8'h00;
RAM[16'h37D7] = 8'h00;
RAM[16'h37D8] = 8'h00;
RAM[16'h37D9] = 8'h00;
RAM[16'h37DA] = 8'h00;
RAM[16'h37DB] = 8'h00;
RAM[16'h37DC] = 8'h00;
RAM[16'h37DD] = 8'h00;
RAM[16'h37DE] = 8'h00;
RAM[16'h37DF] = 8'h00;
RAM[16'h37E0] = 8'h00;
RAM[16'h37E1] = 8'h00;
RAM[16'h37E2] = 8'h00;
RAM[16'h37E3] = 8'h00;
RAM[16'h37E4] = 8'h00;
RAM[16'h37E5] = 8'h00;
RAM[16'h37E6] = 8'h00;
RAM[16'h37E7] = 8'h00;
RAM[16'h37E8] = 8'h00;
RAM[16'h37E9] = 8'h00;
RAM[16'h37EA] = 8'h00;
RAM[16'h37EB] = 8'h00;
RAM[16'h37EC] = 8'h00;
RAM[16'h37ED] = 8'h00;
RAM[16'h37EE] = 8'h00;
RAM[16'h37EF] = 8'h00;
RAM[16'h37F0] = 8'h00;
RAM[16'h37F1] = 8'h00;
RAM[16'h37F2] = 8'h00;
RAM[16'h37F3] = 8'h00;
RAM[16'h37F4] = 8'h00;
RAM[16'h37F5] = 8'h00;
RAM[16'h37F6] = 8'h00;
RAM[16'h37F7] = 8'h00;
RAM[16'h37F8] = 8'h00;
RAM[16'h37F9] = 8'h00;
RAM[16'h37FA] = 8'h00;
RAM[16'h37FB] = 8'h00;
RAM[16'h37FC] = 8'h00;
RAM[16'h37FD] = 8'h00;
RAM[16'h37FE] = 8'h00;
RAM[16'h37FF] = 8'h00;
RAM[16'h3800] = 8'h00;
RAM[16'h3801] = 8'h00;
RAM[16'h3802] = 8'h00;
RAM[16'h3803] = 8'h00;
RAM[16'h3804] = 8'h00;
RAM[16'h3805] = 8'h00;
RAM[16'h3806] = 8'h00;
RAM[16'h3807] = 8'h00;
RAM[16'h3808] = 8'h00;
RAM[16'h3809] = 8'h00;
RAM[16'h380A] = 8'h00;
RAM[16'h380B] = 8'h00;
RAM[16'h380C] = 8'h00;
RAM[16'h380D] = 8'h00;
RAM[16'h380E] = 8'h00;
RAM[16'h380F] = 8'h00;
RAM[16'h3810] = 8'h00;
RAM[16'h3811] = 8'h00;
RAM[16'h3812] = 8'h00;
RAM[16'h3813] = 8'h00;
RAM[16'h3814] = 8'h00;
RAM[16'h3815] = 8'h00;
RAM[16'h3816] = 8'h00;
RAM[16'h3817] = 8'h00;
RAM[16'h3818] = 8'h00;
RAM[16'h3819] = 8'h00;
RAM[16'h381A] = 8'h00;
RAM[16'h381B] = 8'h00;
RAM[16'h381C] = 8'h00;
RAM[16'h381D] = 8'h00;
RAM[16'h381E] = 8'h00;
RAM[16'h381F] = 8'h00;
RAM[16'h3820] = 8'h00;
RAM[16'h3821] = 8'h00;
RAM[16'h3822] = 8'h00;
RAM[16'h3823] = 8'h00;
RAM[16'h3824] = 8'h00;
RAM[16'h3825] = 8'h00;
RAM[16'h3826] = 8'h00;
RAM[16'h3827] = 8'h00;
RAM[16'h3828] = 8'h00;
RAM[16'h3829] = 8'h00;
RAM[16'h382A] = 8'h00;
RAM[16'h382B] = 8'h00;
RAM[16'h382C] = 8'h00;
RAM[16'h382D] = 8'h00;
RAM[16'h382E] = 8'h00;
RAM[16'h382F] = 8'h00;
RAM[16'h3830] = 8'h00;
RAM[16'h3831] = 8'h00;
RAM[16'h3832] = 8'h00;
RAM[16'h3833] = 8'h00;
RAM[16'h3834] = 8'h00;
RAM[16'h3835] = 8'h00;
RAM[16'h3836] = 8'h00;
RAM[16'h3837] = 8'h00;
RAM[16'h3838] = 8'h00;
RAM[16'h3839] = 8'h00;
RAM[16'h383A] = 8'h00;
RAM[16'h383B] = 8'h00;
RAM[16'h383C] = 8'h00;
RAM[16'h383D] = 8'h00;
RAM[16'h383E] = 8'h00;
RAM[16'h383F] = 8'h00;
RAM[16'h3840] = 8'h00;
RAM[16'h3841] = 8'h00;
RAM[16'h3842] = 8'h00;
RAM[16'h3843] = 8'h00;
RAM[16'h3844] = 8'h00;
RAM[16'h3845] = 8'h00;
RAM[16'h3846] = 8'h00;
RAM[16'h3847] = 8'h00;
RAM[16'h3848] = 8'h00;
RAM[16'h3849] = 8'h00;
RAM[16'h384A] = 8'h00;
RAM[16'h384B] = 8'h00;
RAM[16'h384C] = 8'h00;
RAM[16'h384D] = 8'h00;
RAM[16'h384E] = 8'h00;
RAM[16'h384F] = 8'h00;
RAM[16'h3850] = 8'h00;
RAM[16'h3851] = 8'h00;
RAM[16'h3852] = 8'h00;
RAM[16'h3853] = 8'h00;
RAM[16'h3854] = 8'h00;
RAM[16'h3855] = 8'h00;
RAM[16'h3856] = 8'h00;
RAM[16'h3857] = 8'h00;
RAM[16'h3858] = 8'h00;
RAM[16'h3859] = 8'h00;
RAM[16'h385A] = 8'h00;
RAM[16'h385B] = 8'h00;
RAM[16'h385C] = 8'h00;
RAM[16'h385D] = 8'h00;
RAM[16'h385E] = 8'h00;
RAM[16'h385F] = 8'h00;
RAM[16'h3860] = 8'h00;
RAM[16'h3861] = 8'h00;
RAM[16'h3862] = 8'h00;
RAM[16'h3863] = 8'h00;
RAM[16'h3864] = 8'h00;
RAM[16'h3865] = 8'h00;
RAM[16'h3866] = 8'h00;
RAM[16'h3867] = 8'h00;
RAM[16'h3868] = 8'h00;
RAM[16'h3869] = 8'h00;
RAM[16'h386A] = 8'h00;
RAM[16'h386B] = 8'h00;
RAM[16'h386C] = 8'h00;
RAM[16'h386D] = 8'h00;
RAM[16'h386E] = 8'h00;
RAM[16'h386F] = 8'h00;
RAM[16'h3870] = 8'h00;
RAM[16'h3871] = 8'h00;
RAM[16'h3872] = 8'h00;
RAM[16'h3873] = 8'h00;
RAM[16'h3874] = 8'h00;
RAM[16'h3875] = 8'h00;
RAM[16'h3876] = 8'h00;
RAM[16'h3877] = 8'h00;
RAM[16'h3878] = 8'h00;
RAM[16'h3879] = 8'h00;
RAM[16'h387A] = 8'h00;
RAM[16'h387B] = 8'h00;
RAM[16'h387C] = 8'h00;
RAM[16'h387D] = 8'h00;
RAM[16'h387E] = 8'h00;
RAM[16'h387F] = 8'h00;
RAM[16'h3880] = 8'h00;
RAM[16'h3881] = 8'h00;
RAM[16'h3882] = 8'h00;
RAM[16'h3883] = 8'h00;
RAM[16'h3884] = 8'h00;
RAM[16'h3885] = 8'h00;
RAM[16'h3886] = 8'h00;
RAM[16'h3887] = 8'h00;
RAM[16'h3888] = 8'h00;
RAM[16'h3889] = 8'h00;
RAM[16'h388A] = 8'h00;
RAM[16'h388B] = 8'h00;
RAM[16'h388C] = 8'h00;
RAM[16'h388D] = 8'h00;
RAM[16'h388E] = 8'h00;
RAM[16'h388F] = 8'h00;
RAM[16'h3890] = 8'h00;
RAM[16'h3891] = 8'h00;
RAM[16'h3892] = 8'h00;
RAM[16'h3893] = 8'h00;
RAM[16'h3894] = 8'h00;
RAM[16'h3895] = 8'h00;
RAM[16'h3896] = 8'h00;
RAM[16'h3897] = 8'h00;
RAM[16'h3898] = 8'h00;
RAM[16'h3899] = 8'h00;
RAM[16'h389A] = 8'h00;
RAM[16'h389B] = 8'h00;
RAM[16'h389C] = 8'h00;
RAM[16'h389D] = 8'h00;
RAM[16'h389E] = 8'h00;
RAM[16'h389F] = 8'h00;
RAM[16'h38A0] = 8'h00;
RAM[16'h38A1] = 8'h00;
RAM[16'h38A2] = 8'h00;
RAM[16'h38A3] = 8'h00;
RAM[16'h38A4] = 8'h00;
RAM[16'h38A5] = 8'h00;
RAM[16'h38A6] = 8'h00;
RAM[16'h38A7] = 8'h00;
RAM[16'h38A8] = 8'h00;
RAM[16'h38A9] = 8'h00;
RAM[16'h38AA] = 8'h00;
RAM[16'h38AB] = 8'h00;
RAM[16'h38AC] = 8'h00;
RAM[16'h38AD] = 8'h00;
RAM[16'h38AE] = 8'h00;
RAM[16'h38AF] = 8'h00;
RAM[16'h38B0] = 8'h00;
RAM[16'h38B1] = 8'h00;
RAM[16'h38B2] = 8'h00;
RAM[16'h38B3] = 8'h00;
RAM[16'h38B4] = 8'h00;
RAM[16'h38B5] = 8'h00;
RAM[16'h38B6] = 8'h00;
RAM[16'h38B7] = 8'h00;
RAM[16'h38B8] = 8'h00;
RAM[16'h38B9] = 8'h00;
RAM[16'h38BA] = 8'h00;
RAM[16'h38BB] = 8'h00;
RAM[16'h38BC] = 8'h00;
RAM[16'h38BD] = 8'h00;
RAM[16'h38BE] = 8'h00;
RAM[16'h38BF] = 8'h00;
RAM[16'h38C0] = 8'h00;
RAM[16'h38C1] = 8'h00;
RAM[16'h38C2] = 8'h00;
RAM[16'h38C3] = 8'h00;
RAM[16'h38C4] = 8'h00;
RAM[16'h38C5] = 8'h00;
RAM[16'h38C6] = 8'h00;
RAM[16'h38C7] = 8'h00;
RAM[16'h38C8] = 8'h00;
RAM[16'h38C9] = 8'h00;
RAM[16'h38CA] = 8'h00;
RAM[16'h38CB] = 8'h00;
RAM[16'h38CC] = 8'h00;
RAM[16'h38CD] = 8'h00;
RAM[16'h38CE] = 8'h00;
RAM[16'h38CF] = 8'h00;
RAM[16'h38D0] = 8'h00;
RAM[16'h38D1] = 8'h00;
RAM[16'h38D2] = 8'h00;
RAM[16'h38D3] = 8'h00;
RAM[16'h38D4] = 8'h00;
RAM[16'h38D5] = 8'h00;
RAM[16'h38D6] = 8'h00;
RAM[16'h38D7] = 8'h00;
RAM[16'h38D8] = 8'h00;
RAM[16'h38D9] = 8'h00;
RAM[16'h38DA] = 8'h00;
RAM[16'h38DB] = 8'h00;
RAM[16'h38DC] = 8'h00;
RAM[16'h38DD] = 8'h00;
RAM[16'h38DE] = 8'h00;
RAM[16'h38DF] = 8'h00;
RAM[16'h38E0] = 8'h00;
RAM[16'h38E1] = 8'h00;
RAM[16'h38E2] = 8'h00;
RAM[16'h38E3] = 8'h00;
RAM[16'h38E4] = 8'h00;
RAM[16'h38E5] = 8'h00;
RAM[16'h38E6] = 8'h00;
RAM[16'h38E7] = 8'h00;
RAM[16'h38E8] = 8'h00;
RAM[16'h38E9] = 8'h00;
RAM[16'h38EA] = 8'h00;
RAM[16'h38EB] = 8'h00;
RAM[16'h38EC] = 8'h00;
RAM[16'h38ED] = 8'h00;
RAM[16'h38EE] = 8'h00;
RAM[16'h38EF] = 8'h00;
RAM[16'h38F0] = 8'h00;
RAM[16'h38F1] = 8'h00;
RAM[16'h38F2] = 8'h00;
RAM[16'h38F3] = 8'h00;
RAM[16'h38F4] = 8'h00;
RAM[16'h38F5] = 8'h00;
RAM[16'h38F6] = 8'h00;
RAM[16'h38F7] = 8'h00;
RAM[16'h38F8] = 8'h00;
RAM[16'h38F9] = 8'h00;
RAM[16'h38FA] = 8'h00;
RAM[16'h38FB] = 8'h00;
RAM[16'h38FC] = 8'h00;
RAM[16'h38FD] = 8'h00;
RAM[16'h38FE] = 8'h00;
RAM[16'h38FF] = 8'h00;
RAM[16'h3900] = 8'h00;
RAM[16'h3901] = 8'h00;
RAM[16'h3902] = 8'h00;
RAM[16'h3903] = 8'h00;
RAM[16'h3904] = 8'h00;
RAM[16'h3905] = 8'h00;
RAM[16'h3906] = 8'h00;
RAM[16'h3907] = 8'h00;
RAM[16'h3908] = 8'h00;
RAM[16'h3909] = 8'h00;
RAM[16'h390A] = 8'h00;
RAM[16'h390B] = 8'h00;
RAM[16'h390C] = 8'h00;
RAM[16'h390D] = 8'h00;
RAM[16'h390E] = 8'h00;
RAM[16'h390F] = 8'h00;
RAM[16'h3910] = 8'h00;
RAM[16'h3911] = 8'h00;
RAM[16'h3912] = 8'h00;
RAM[16'h3913] = 8'h00;
RAM[16'h3914] = 8'h00;
RAM[16'h3915] = 8'h00;
RAM[16'h3916] = 8'h00;
RAM[16'h3917] = 8'h00;
RAM[16'h3918] = 8'h00;
RAM[16'h3919] = 8'h00;
RAM[16'h391A] = 8'h00;
RAM[16'h391B] = 8'h00;
RAM[16'h391C] = 8'h00;
RAM[16'h391D] = 8'h00;
RAM[16'h391E] = 8'h00;
RAM[16'h391F] = 8'h00;
RAM[16'h3920] = 8'h00;
RAM[16'h3921] = 8'h00;
RAM[16'h3922] = 8'h00;
RAM[16'h3923] = 8'h00;
RAM[16'h3924] = 8'h00;
RAM[16'h3925] = 8'h00;
RAM[16'h3926] = 8'h00;
RAM[16'h3927] = 8'h00;
RAM[16'h3928] = 8'h00;
RAM[16'h3929] = 8'h00;
RAM[16'h392A] = 8'h00;
RAM[16'h392B] = 8'h00;
RAM[16'h392C] = 8'h00;
RAM[16'h392D] = 8'h00;
RAM[16'h392E] = 8'h00;
RAM[16'h392F] = 8'h00;
RAM[16'h3930] = 8'h00;
RAM[16'h3931] = 8'h00;
RAM[16'h3932] = 8'h00;
RAM[16'h3933] = 8'h00;
RAM[16'h3934] = 8'h00;
RAM[16'h3935] = 8'h00;
RAM[16'h3936] = 8'h00;
RAM[16'h3937] = 8'h00;
RAM[16'h3938] = 8'h00;
RAM[16'h3939] = 8'h00;
RAM[16'h393A] = 8'h00;
RAM[16'h393B] = 8'h00;
RAM[16'h393C] = 8'h00;
RAM[16'h393D] = 8'h00;
RAM[16'h393E] = 8'h00;
RAM[16'h393F] = 8'h00;
RAM[16'h3940] = 8'h00;
RAM[16'h3941] = 8'h00;
RAM[16'h3942] = 8'h00;
RAM[16'h3943] = 8'h00;
RAM[16'h3944] = 8'h00;
RAM[16'h3945] = 8'h00;
RAM[16'h3946] = 8'h00;
RAM[16'h3947] = 8'h00;
RAM[16'h3948] = 8'h00;
RAM[16'h3949] = 8'h00;
RAM[16'h394A] = 8'h00;
RAM[16'h394B] = 8'h00;
RAM[16'h394C] = 8'h00;
RAM[16'h394D] = 8'h00;
RAM[16'h394E] = 8'h00;
RAM[16'h394F] = 8'h00;
RAM[16'h3950] = 8'h00;
RAM[16'h3951] = 8'h00;
RAM[16'h3952] = 8'h00;
RAM[16'h3953] = 8'h00;
RAM[16'h3954] = 8'h00;
RAM[16'h3955] = 8'h00;
RAM[16'h3956] = 8'h00;
RAM[16'h3957] = 8'h00;
RAM[16'h3958] = 8'h00;
RAM[16'h3959] = 8'h00;
RAM[16'h395A] = 8'h00;
RAM[16'h395B] = 8'h00;
RAM[16'h395C] = 8'h00;
RAM[16'h395D] = 8'h00;
RAM[16'h395E] = 8'h00;
RAM[16'h395F] = 8'h00;
RAM[16'h3960] = 8'h00;
RAM[16'h3961] = 8'h00;
RAM[16'h3962] = 8'h00;
RAM[16'h3963] = 8'h00;
RAM[16'h3964] = 8'h00;
RAM[16'h3965] = 8'h00;
RAM[16'h3966] = 8'h00;
RAM[16'h3967] = 8'h00;
RAM[16'h3968] = 8'h00;
RAM[16'h3969] = 8'h00;
RAM[16'h396A] = 8'h00;
RAM[16'h396B] = 8'h00;
RAM[16'h396C] = 8'h00;
RAM[16'h396D] = 8'h00;
RAM[16'h396E] = 8'h00;
RAM[16'h396F] = 8'h00;
RAM[16'h3970] = 8'h00;
RAM[16'h3971] = 8'h00;
RAM[16'h3972] = 8'h00;
RAM[16'h3973] = 8'h00;
RAM[16'h3974] = 8'h00;
RAM[16'h3975] = 8'h00;
RAM[16'h3976] = 8'h00;
RAM[16'h3977] = 8'h00;
RAM[16'h3978] = 8'h00;
RAM[16'h3979] = 8'h00;
RAM[16'h397A] = 8'h00;
RAM[16'h397B] = 8'h00;
RAM[16'h397C] = 8'h00;
RAM[16'h397D] = 8'h00;
RAM[16'h397E] = 8'h00;
RAM[16'h397F] = 8'h00;
RAM[16'h3980] = 8'h00;
RAM[16'h3981] = 8'h00;
RAM[16'h3982] = 8'h00;
RAM[16'h3983] = 8'h00;
RAM[16'h3984] = 8'h00;
RAM[16'h3985] = 8'h00;
RAM[16'h3986] = 8'h00;
RAM[16'h3987] = 8'h00;
RAM[16'h3988] = 8'h00;
RAM[16'h3989] = 8'h00;
RAM[16'h398A] = 8'h00;
RAM[16'h398B] = 8'h00;
RAM[16'h398C] = 8'h00;
RAM[16'h398D] = 8'h00;
RAM[16'h398E] = 8'h00;
RAM[16'h398F] = 8'h00;
RAM[16'h3990] = 8'h00;
RAM[16'h3991] = 8'h00;
RAM[16'h3992] = 8'h00;
RAM[16'h3993] = 8'h00;
RAM[16'h3994] = 8'h00;
RAM[16'h3995] = 8'h00;
RAM[16'h3996] = 8'h00;
RAM[16'h3997] = 8'h00;
RAM[16'h3998] = 8'h00;
RAM[16'h3999] = 8'h00;
RAM[16'h399A] = 8'h00;
RAM[16'h399B] = 8'h00;
RAM[16'h399C] = 8'h00;
RAM[16'h399D] = 8'h00;
RAM[16'h399E] = 8'h00;
RAM[16'h399F] = 8'h00;
RAM[16'h39A0] = 8'h00;
RAM[16'h39A1] = 8'h00;
RAM[16'h39A2] = 8'h00;
RAM[16'h39A3] = 8'h00;
RAM[16'h39A4] = 8'h00;
RAM[16'h39A5] = 8'h00;
RAM[16'h39A6] = 8'h00;
RAM[16'h39A7] = 8'h00;
RAM[16'h39A8] = 8'h00;
RAM[16'h39A9] = 8'h00;
RAM[16'h39AA] = 8'h00;
RAM[16'h39AB] = 8'h00;
RAM[16'h39AC] = 8'h00;
RAM[16'h39AD] = 8'h00;
RAM[16'h39AE] = 8'h00;
RAM[16'h39AF] = 8'h00;
RAM[16'h39B0] = 8'h00;
RAM[16'h39B1] = 8'h00;
RAM[16'h39B2] = 8'h00;
RAM[16'h39B3] = 8'h00;
RAM[16'h39B4] = 8'h00;
RAM[16'h39B5] = 8'h00;
RAM[16'h39B6] = 8'h00;
RAM[16'h39B7] = 8'h00;
RAM[16'h39B8] = 8'h00;
RAM[16'h39B9] = 8'h00;
RAM[16'h39BA] = 8'h00;
RAM[16'h39BB] = 8'h00;
RAM[16'h39BC] = 8'h00;
RAM[16'h39BD] = 8'h00;
RAM[16'h39BE] = 8'h00;
RAM[16'h39BF] = 8'h00;
RAM[16'h39C0] = 8'h00;
RAM[16'h39C1] = 8'h00;
RAM[16'h39C2] = 8'h00;
RAM[16'h39C3] = 8'h00;
RAM[16'h39C4] = 8'h00;
RAM[16'h39C5] = 8'h00;
RAM[16'h39C6] = 8'h00;
RAM[16'h39C7] = 8'h00;
RAM[16'h39C8] = 8'h00;
RAM[16'h39C9] = 8'h00;
RAM[16'h39CA] = 8'h00;
RAM[16'h39CB] = 8'h00;
RAM[16'h39CC] = 8'h00;
RAM[16'h39CD] = 8'h00;
RAM[16'h39CE] = 8'h00;
RAM[16'h39CF] = 8'h00;
RAM[16'h39D0] = 8'h00;
RAM[16'h39D1] = 8'h00;
RAM[16'h39D2] = 8'h00;
RAM[16'h39D3] = 8'h00;
RAM[16'h39D4] = 8'h00;
RAM[16'h39D5] = 8'h00;
RAM[16'h39D6] = 8'h00;
RAM[16'h39D7] = 8'h00;
RAM[16'h39D8] = 8'h00;
RAM[16'h39D9] = 8'h00;
RAM[16'h39DA] = 8'h00;
RAM[16'h39DB] = 8'h00;
RAM[16'h39DC] = 8'h00;
RAM[16'h39DD] = 8'h00;
RAM[16'h39DE] = 8'h00;
RAM[16'h39DF] = 8'h00;
RAM[16'h39E0] = 8'h00;
RAM[16'h39E1] = 8'h00;
RAM[16'h39E2] = 8'h00;
RAM[16'h39E3] = 8'h00;
RAM[16'h39E4] = 8'h00;
RAM[16'h39E5] = 8'h00;
RAM[16'h39E6] = 8'h00;
RAM[16'h39E7] = 8'h00;
RAM[16'h39E8] = 8'h00;
RAM[16'h39E9] = 8'h00;
RAM[16'h39EA] = 8'h00;
RAM[16'h39EB] = 8'h00;
RAM[16'h39EC] = 8'h00;
RAM[16'h39ED] = 8'h00;
RAM[16'h39EE] = 8'h00;
RAM[16'h39EF] = 8'h00;
RAM[16'h39F0] = 8'h00;
RAM[16'h39F1] = 8'h00;
RAM[16'h39F2] = 8'h00;
RAM[16'h39F3] = 8'h00;
RAM[16'h39F4] = 8'h00;
RAM[16'h39F5] = 8'h00;
RAM[16'h39F6] = 8'h00;
RAM[16'h39F7] = 8'h00;
RAM[16'h39F8] = 8'h00;
RAM[16'h39F9] = 8'h00;
RAM[16'h39FA] = 8'h00;
RAM[16'h39FB] = 8'h00;
RAM[16'h39FC] = 8'h00;
RAM[16'h39FD] = 8'h00;
RAM[16'h39FE] = 8'h00;
RAM[16'h39FF] = 8'h00;
RAM[16'h3A00] = 8'h00;
RAM[16'h3A01] = 8'h00;
RAM[16'h3A02] = 8'h00;
RAM[16'h3A03] = 8'h00;
RAM[16'h3A04] = 8'h00;
RAM[16'h3A05] = 8'h00;
RAM[16'h3A06] = 8'h00;
RAM[16'h3A07] = 8'h00;
RAM[16'h3A08] = 8'h00;
RAM[16'h3A09] = 8'h00;
RAM[16'h3A0A] = 8'h00;
RAM[16'h3A0B] = 8'h00;
RAM[16'h3A0C] = 8'h00;
RAM[16'h3A0D] = 8'h00;
RAM[16'h3A0E] = 8'h00;
RAM[16'h3A0F] = 8'h00;
RAM[16'h3A10] = 8'h00;
RAM[16'h3A11] = 8'h00;
RAM[16'h3A12] = 8'h00;
RAM[16'h3A13] = 8'h00;
RAM[16'h3A14] = 8'h00;
RAM[16'h3A15] = 8'h00;
RAM[16'h3A16] = 8'h00;
RAM[16'h3A17] = 8'h00;
RAM[16'h3A18] = 8'h00;
RAM[16'h3A19] = 8'h00;
RAM[16'h3A1A] = 8'h00;
RAM[16'h3A1B] = 8'h00;
RAM[16'h3A1C] = 8'h00;
RAM[16'h3A1D] = 8'h00;
RAM[16'h3A1E] = 8'h00;
RAM[16'h3A1F] = 8'h00;
RAM[16'h3A20] = 8'h00;
RAM[16'h3A21] = 8'h00;
RAM[16'h3A22] = 8'h00;
RAM[16'h3A23] = 8'h00;
RAM[16'h3A24] = 8'h00;
RAM[16'h3A25] = 8'h00;
RAM[16'h3A26] = 8'h00;
RAM[16'h3A27] = 8'h00;
RAM[16'h3A28] = 8'h00;
RAM[16'h3A29] = 8'h00;
RAM[16'h3A2A] = 8'h00;
RAM[16'h3A2B] = 8'h00;
RAM[16'h3A2C] = 8'h00;
RAM[16'h3A2D] = 8'h00;
RAM[16'h3A2E] = 8'h00;
RAM[16'h3A2F] = 8'h00;
RAM[16'h3A30] = 8'h00;
RAM[16'h3A31] = 8'h00;
RAM[16'h3A32] = 8'h00;
RAM[16'h3A33] = 8'h00;
RAM[16'h3A34] = 8'h00;
RAM[16'h3A35] = 8'h00;
RAM[16'h3A36] = 8'h00;
RAM[16'h3A37] = 8'h00;
RAM[16'h3A38] = 8'h00;
RAM[16'h3A39] = 8'h00;
RAM[16'h3A3A] = 8'h00;
RAM[16'h3A3B] = 8'h00;
RAM[16'h3A3C] = 8'h00;
RAM[16'h3A3D] = 8'h00;
RAM[16'h3A3E] = 8'h00;
RAM[16'h3A3F] = 8'h00;
RAM[16'h3A40] = 8'h00;
RAM[16'h3A41] = 8'h00;
RAM[16'h3A42] = 8'h00;
RAM[16'h3A43] = 8'h00;
RAM[16'h3A44] = 8'h00;
RAM[16'h3A45] = 8'h00;
RAM[16'h3A46] = 8'h00;
RAM[16'h3A47] = 8'h00;
RAM[16'h3A48] = 8'h00;
RAM[16'h3A49] = 8'h00;
RAM[16'h3A4A] = 8'h00;
RAM[16'h3A4B] = 8'h00;
RAM[16'h3A4C] = 8'h00;
RAM[16'h3A4D] = 8'h00;
RAM[16'h3A4E] = 8'h00;
RAM[16'h3A4F] = 8'h00;
RAM[16'h3A50] = 8'h00;
RAM[16'h3A51] = 8'h00;
RAM[16'h3A52] = 8'h00;
RAM[16'h3A53] = 8'h00;
RAM[16'h3A54] = 8'h00;
RAM[16'h3A55] = 8'h00;
RAM[16'h3A56] = 8'h00;
RAM[16'h3A57] = 8'h00;
RAM[16'h3A58] = 8'h00;
RAM[16'h3A59] = 8'h00;
RAM[16'h3A5A] = 8'h00;
RAM[16'h3A5B] = 8'h00;
RAM[16'h3A5C] = 8'h00;
RAM[16'h3A5D] = 8'h00;
RAM[16'h3A5E] = 8'h00;
RAM[16'h3A5F] = 8'h00;
RAM[16'h3A60] = 8'h00;
RAM[16'h3A61] = 8'h00;
RAM[16'h3A62] = 8'h00;
RAM[16'h3A63] = 8'h00;
RAM[16'h3A64] = 8'h00;
RAM[16'h3A65] = 8'h00;
RAM[16'h3A66] = 8'h00;
RAM[16'h3A67] = 8'h00;
RAM[16'h3A68] = 8'h00;
RAM[16'h3A69] = 8'h00;
RAM[16'h3A6A] = 8'h00;
RAM[16'h3A6B] = 8'h00;
RAM[16'h3A6C] = 8'h00;
RAM[16'h3A6D] = 8'h00;
RAM[16'h3A6E] = 8'h00;
RAM[16'h3A6F] = 8'h00;
RAM[16'h3A70] = 8'h00;
RAM[16'h3A71] = 8'h00;
RAM[16'h3A72] = 8'h00;
RAM[16'h3A73] = 8'h00;
RAM[16'h3A74] = 8'h00;
RAM[16'h3A75] = 8'h00;
RAM[16'h3A76] = 8'h00;
RAM[16'h3A77] = 8'h00;
RAM[16'h3A78] = 8'h00;
RAM[16'h3A79] = 8'h00;
RAM[16'h3A7A] = 8'h00;
RAM[16'h3A7B] = 8'h00;
RAM[16'h3A7C] = 8'h00;
RAM[16'h3A7D] = 8'h00;
RAM[16'h3A7E] = 8'h00;
RAM[16'h3A7F] = 8'h00;
RAM[16'h3A80] = 8'h00;
RAM[16'h3A81] = 8'h00;
RAM[16'h3A82] = 8'h00;
RAM[16'h3A83] = 8'h00;
RAM[16'h3A84] = 8'h00;
RAM[16'h3A85] = 8'h00;
RAM[16'h3A86] = 8'h00;
RAM[16'h3A87] = 8'h00;
RAM[16'h3A88] = 8'h00;
RAM[16'h3A89] = 8'h00;
RAM[16'h3A8A] = 8'h00;
RAM[16'h3A8B] = 8'h00;
RAM[16'h3A8C] = 8'h00;
RAM[16'h3A8D] = 8'h00;
RAM[16'h3A8E] = 8'h00;
RAM[16'h3A8F] = 8'h00;
RAM[16'h3A90] = 8'h00;
RAM[16'h3A91] = 8'h00;
RAM[16'h3A92] = 8'h00;
RAM[16'h3A93] = 8'h00;
RAM[16'h3A94] = 8'h00;
RAM[16'h3A95] = 8'h00;
RAM[16'h3A96] = 8'h00;
RAM[16'h3A97] = 8'h00;
RAM[16'h3A98] = 8'h00;
RAM[16'h3A99] = 8'h00;
RAM[16'h3A9A] = 8'h00;
RAM[16'h3A9B] = 8'h00;
RAM[16'h3A9C] = 8'h00;
RAM[16'h3A9D] = 8'h00;
RAM[16'h3A9E] = 8'h00;
RAM[16'h3A9F] = 8'h00;
RAM[16'h3AA0] = 8'h00;
RAM[16'h3AA1] = 8'h00;
RAM[16'h3AA2] = 8'h00;
RAM[16'h3AA3] = 8'h00;
RAM[16'h3AA4] = 8'h00;
RAM[16'h3AA5] = 8'h00;
RAM[16'h3AA6] = 8'h00;
RAM[16'h3AA7] = 8'h00;
RAM[16'h3AA8] = 8'h00;
RAM[16'h3AA9] = 8'h00;
RAM[16'h3AAA] = 8'h00;
RAM[16'h3AAB] = 8'h00;
RAM[16'h3AAC] = 8'h00;
RAM[16'h3AAD] = 8'h00;
RAM[16'h3AAE] = 8'h00;
RAM[16'h3AAF] = 8'h00;
RAM[16'h3AB0] = 8'h00;
RAM[16'h3AB1] = 8'h00;
RAM[16'h3AB2] = 8'h00;
RAM[16'h3AB3] = 8'h00;
RAM[16'h3AB4] = 8'h00;
RAM[16'h3AB5] = 8'h00;
RAM[16'h3AB6] = 8'h00;
RAM[16'h3AB7] = 8'h00;
RAM[16'h3AB8] = 8'h00;
RAM[16'h3AB9] = 8'h00;
RAM[16'h3ABA] = 8'h00;
RAM[16'h3ABB] = 8'h00;
RAM[16'h3ABC] = 8'h00;
RAM[16'h3ABD] = 8'h00;
RAM[16'h3ABE] = 8'h00;
RAM[16'h3ABF] = 8'h00;
RAM[16'h3AC0] = 8'h00;
RAM[16'h3AC1] = 8'h00;
RAM[16'h3AC2] = 8'h00;
RAM[16'h3AC3] = 8'h00;
RAM[16'h3AC4] = 8'h00;
RAM[16'h3AC5] = 8'h00;
RAM[16'h3AC6] = 8'h00;
RAM[16'h3AC7] = 8'h00;
RAM[16'h3AC8] = 8'h00;
RAM[16'h3AC9] = 8'h00;
RAM[16'h3ACA] = 8'h00;
RAM[16'h3ACB] = 8'h00;
RAM[16'h3ACC] = 8'h00;
RAM[16'h3ACD] = 8'h00;
RAM[16'h3ACE] = 8'h00;
RAM[16'h3ACF] = 8'h00;
RAM[16'h3AD0] = 8'h00;
RAM[16'h3AD1] = 8'h00;
RAM[16'h3AD2] = 8'h00;
RAM[16'h3AD3] = 8'h00;
RAM[16'h3AD4] = 8'h00;
RAM[16'h3AD5] = 8'h00;
RAM[16'h3AD6] = 8'h00;
RAM[16'h3AD7] = 8'h00;
RAM[16'h3AD8] = 8'h00;
RAM[16'h3AD9] = 8'h00;
RAM[16'h3ADA] = 8'h00;
RAM[16'h3ADB] = 8'h00;
RAM[16'h3ADC] = 8'h00;
RAM[16'h3ADD] = 8'h00;
RAM[16'h3ADE] = 8'h00;
RAM[16'h3ADF] = 8'h00;
RAM[16'h3AE0] = 8'h00;
RAM[16'h3AE1] = 8'h00;
RAM[16'h3AE2] = 8'h00;
RAM[16'h3AE3] = 8'h00;
RAM[16'h3AE4] = 8'h00;
RAM[16'h3AE5] = 8'h00;
RAM[16'h3AE6] = 8'h00;
RAM[16'h3AE7] = 8'h00;
RAM[16'h3AE8] = 8'h00;
RAM[16'h3AE9] = 8'h00;
RAM[16'h3AEA] = 8'h00;
RAM[16'h3AEB] = 8'h00;
RAM[16'h3AEC] = 8'h00;
RAM[16'h3AED] = 8'h00;
RAM[16'h3AEE] = 8'h00;
RAM[16'h3AEF] = 8'h00;
RAM[16'h3AF0] = 8'h00;
RAM[16'h3AF1] = 8'h00;
RAM[16'h3AF2] = 8'h00;
RAM[16'h3AF3] = 8'h00;
RAM[16'h3AF4] = 8'h00;
RAM[16'h3AF5] = 8'h00;
RAM[16'h3AF6] = 8'h00;
RAM[16'h3AF7] = 8'h00;
RAM[16'h3AF8] = 8'h00;
RAM[16'h3AF9] = 8'h00;
RAM[16'h3AFA] = 8'h00;
RAM[16'h3AFB] = 8'h00;
RAM[16'h3AFC] = 8'h00;
RAM[16'h3AFD] = 8'h00;
RAM[16'h3AFE] = 8'h00;
RAM[16'h3AFF] = 8'h00;
RAM[16'h3B00] = 8'h00;
RAM[16'h3B01] = 8'h00;
RAM[16'h3B02] = 8'h00;
RAM[16'h3B03] = 8'h00;
RAM[16'h3B04] = 8'h00;
RAM[16'h3B05] = 8'h00;
RAM[16'h3B06] = 8'h00;
RAM[16'h3B07] = 8'h00;
RAM[16'h3B08] = 8'h00;
RAM[16'h3B09] = 8'h00;
RAM[16'h3B0A] = 8'h00;
RAM[16'h3B0B] = 8'h00;
RAM[16'h3B0C] = 8'h00;
RAM[16'h3B0D] = 8'h00;
RAM[16'h3B0E] = 8'h00;
RAM[16'h3B0F] = 8'h00;
RAM[16'h3B10] = 8'h00;
RAM[16'h3B11] = 8'h00;
RAM[16'h3B12] = 8'h00;
RAM[16'h3B13] = 8'h00;
RAM[16'h3B14] = 8'h00;
RAM[16'h3B15] = 8'h00;
RAM[16'h3B16] = 8'h00;
RAM[16'h3B17] = 8'h00;
RAM[16'h3B18] = 8'h00;
RAM[16'h3B19] = 8'h00;
RAM[16'h3B1A] = 8'h00;
RAM[16'h3B1B] = 8'h00;
RAM[16'h3B1C] = 8'h00;
RAM[16'h3B1D] = 8'h00;
RAM[16'h3B1E] = 8'h00;
RAM[16'h3B1F] = 8'h00;
RAM[16'h3B20] = 8'h00;
RAM[16'h3B21] = 8'h00;
RAM[16'h3B22] = 8'h00;
RAM[16'h3B23] = 8'h00;
RAM[16'h3B24] = 8'h00;
RAM[16'h3B25] = 8'h00;
RAM[16'h3B26] = 8'h00;
RAM[16'h3B27] = 8'h00;
RAM[16'h3B28] = 8'h00;
RAM[16'h3B29] = 8'h00;
RAM[16'h3B2A] = 8'h00;
RAM[16'h3B2B] = 8'h00;
RAM[16'h3B2C] = 8'h00;
RAM[16'h3B2D] = 8'h00;
RAM[16'h3B2E] = 8'h00;
RAM[16'h3B2F] = 8'h00;
RAM[16'h3B30] = 8'h00;
RAM[16'h3B31] = 8'h00;
RAM[16'h3B32] = 8'h00;
RAM[16'h3B33] = 8'h00;
RAM[16'h3B34] = 8'h00;
RAM[16'h3B35] = 8'h00;
RAM[16'h3B36] = 8'h00;
RAM[16'h3B37] = 8'h00;
RAM[16'h3B38] = 8'h00;
RAM[16'h3B39] = 8'h00;
RAM[16'h3B3A] = 8'h00;
RAM[16'h3B3B] = 8'h00;
RAM[16'h3B3C] = 8'h00;
RAM[16'h3B3D] = 8'h00;
RAM[16'h3B3E] = 8'h00;
RAM[16'h3B3F] = 8'h00;
RAM[16'h3B40] = 8'h00;
RAM[16'h3B41] = 8'h00;
RAM[16'h3B42] = 8'h00;
RAM[16'h3B43] = 8'h00;
RAM[16'h3B44] = 8'h00;
RAM[16'h3B45] = 8'h00;
RAM[16'h3B46] = 8'h00;
RAM[16'h3B47] = 8'h00;
RAM[16'h3B48] = 8'h00;
RAM[16'h3B49] = 8'h00;
RAM[16'h3B4A] = 8'h00;
RAM[16'h3B4B] = 8'h00;
RAM[16'h3B4C] = 8'h00;
RAM[16'h3B4D] = 8'h00;
RAM[16'h3B4E] = 8'h00;
RAM[16'h3B4F] = 8'h00;
RAM[16'h3B50] = 8'h00;
RAM[16'h3B51] = 8'h00;
RAM[16'h3B52] = 8'h00;
RAM[16'h3B53] = 8'h00;
RAM[16'h3B54] = 8'h00;
RAM[16'h3B55] = 8'h00;
RAM[16'h3B56] = 8'h00;
RAM[16'h3B57] = 8'h00;
RAM[16'h3B58] = 8'h00;
RAM[16'h3B59] = 8'h00;
RAM[16'h3B5A] = 8'h00;
RAM[16'h3B5B] = 8'h00;
RAM[16'h3B5C] = 8'h00;
RAM[16'h3B5D] = 8'h00;
RAM[16'h3B5E] = 8'h00;
RAM[16'h3B5F] = 8'h00;
RAM[16'h3B60] = 8'h00;
RAM[16'h3B61] = 8'h00;
RAM[16'h3B62] = 8'h00;
RAM[16'h3B63] = 8'h00;
RAM[16'h3B64] = 8'h00;
RAM[16'h3B65] = 8'h00;
RAM[16'h3B66] = 8'h00;
RAM[16'h3B67] = 8'h00;
RAM[16'h3B68] = 8'h00;
RAM[16'h3B69] = 8'h00;
RAM[16'h3B6A] = 8'h00;
RAM[16'h3B6B] = 8'h00;
RAM[16'h3B6C] = 8'h00;
RAM[16'h3B6D] = 8'h00;
RAM[16'h3B6E] = 8'h00;
RAM[16'h3B6F] = 8'h00;
RAM[16'h3B70] = 8'h00;
RAM[16'h3B71] = 8'h00;
RAM[16'h3B72] = 8'h00;
RAM[16'h3B73] = 8'h00;
RAM[16'h3B74] = 8'h00;
RAM[16'h3B75] = 8'h00;
RAM[16'h3B76] = 8'h00;
RAM[16'h3B77] = 8'h00;
RAM[16'h3B78] = 8'h00;
RAM[16'h3B79] = 8'h00;
RAM[16'h3B7A] = 8'h00;
RAM[16'h3B7B] = 8'h00;
RAM[16'h3B7C] = 8'h00;
RAM[16'h3B7D] = 8'h00;
RAM[16'h3B7E] = 8'h00;
RAM[16'h3B7F] = 8'h00;
RAM[16'h3B80] = 8'h00;
RAM[16'h3B81] = 8'h00;
RAM[16'h3B82] = 8'h00;
RAM[16'h3B83] = 8'h00;
RAM[16'h3B84] = 8'h00;
RAM[16'h3B85] = 8'h00;
RAM[16'h3B86] = 8'h00;
RAM[16'h3B87] = 8'h00;
RAM[16'h3B88] = 8'h00;
RAM[16'h3B89] = 8'h00;
RAM[16'h3B8A] = 8'h00;
RAM[16'h3B8B] = 8'h00;
RAM[16'h3B8C] = 8'h00;
RAM[16'h3B8D] = 8'h00;
RAM[16'h3B8E] = 8'h00;
RAM[16'h3B8F] = 8'h00;
RAM[16'h3B90] = 8'h00;
RAM[16'h3B91] = 8'h00;
RAM[16'h3B92] = 8'h00;
RAM[16'h3B93] = 8'h00;
RAM[16'h3B94] = 8'h00;
RAM[16'h3B95] = 8'h00;
RAM[16'h3B96] = 8'h00;
RAM[16'h3B97] = 8'h00;
RAM[16'h3B98] = 8'h00;
RAM[16'h3B99] = 8'h00;
RAM[16'h3B9A] = 8'h00;
RAM[16'h3B9B] = 8'h00;
RAM[16'h3B9C] = 8'h00;
RAM[16'h3B9D] = 8'h00;
RAM[16'h3B9E] = 8'h00;
RAM[16'h3B9F] = 8'h00;
RAM[16'h3BA0] = 8'h00;
RAM[16'h3BA1] = 8'h00;
RAM[16'h3BA2] = 8'h00;
RAM[16'h3BA3] = 8'h00;
RAM[16'h3BA4] = 8'h00;
RAM[16'h3BA5] = 8'h00;
RAM[16'h3BA6] = 8'h00;
RAM[16'h3BA7] = 8'h00;
RAM[16'h3BA8] = 8'h00;
RAM[16'h3BA9] = 8'h00;
RAM[16'h3BAA] = 8'h00;
RAM[16'h3BAB] = 8'h00;
RAM[16'h3BAC] = 8'h00;
RAM[16'h3BAD] = 8'h00;
RAM[16'h3BAE] = 8'h00;
RAM[16'h3BAF] = 8'h00;
RAM[16'h3BB0] = 8'h00;
RAM[16'h3BB1] = 8'h00;
RAM[16'h3BB2] = 8'h00;
RAM[16'h3BB3] = 8'h00;
RAM[16'h3BB4] = 8'h00;
RAM[16'h3BB5] = 8'h00;
RAM[16'h3BB6] = 8'h00;
RAM[16'h3BB7] = 8'h00;
RAM[16'h3BB8] = 8'h00;
RAM[16'h3BB9] = 8'h00;
RAM[16'h3BBA] = 8'h00;
RAM[16'h3BBB] = 8'h00;
RAM[16'h3BBC] = 8'h00;
RAM[16'h3BBD] = 8'h00;
RAM[16'h3BBE] = 8'h00;
RAM[16'h3BBF] = 8'h00;
RAM[16'h3BC0] = 8'h00;
RAM[16'h3BC1] = 8'h00;
RAM[16'h3BC2] = 8'h00;
RAM[16'h3BC3] = 8'h00;
RAM[16'h3BC4] = 8'h00;
RAM[16'h3BC5] = 8'h00;
RAM[16'h3BC6] = 8'h00;
RAM[16'h3BC7] = 8'h00;
RAM[16'h3BC8] = 8'h00;
RAM[16'h3BC9] = 8'h00;
RAM[16'h3BCA] = 8'h00;
RAM[16'h3BCB] = 8'h00;
RAM[16'h3BCC] = 8'h00;
RAM[16'h3BCD] = 8'h00;
RAM[16'h3BCE] = 8'h00;
RAM[16'h3BCF] = 8'h00;
RAM[16'h3BD0] = 8'h00;
RAM[16'h3BD1] = 8'h00;
RAM[16'h3BD2] = 8'h00;
RAM[16'h3BD3] = 8'h00;
RAM[16'h3BD4] = 8'h00;
RAM[16'h3BD5] = 8'h00;
RAM[16'h3BD6] = 8'h00;
RAM[16'h3BD7] = 8'h00;
RAM[16'h3BD8] = 8'h00;
RAM[16'h3BD9] = 8'h00;
RAM[16'h3BDA] = 8'h00;
RAM[16'h3BDB] = 8'h00;
RAM[16'h3BDC] = 8'h00;
RAM[16'h3BDD] = 8'h00;
RAM[16'h3BDE] = 8'h00;
RAM[16'h3BDF] = 8'h00;
RAM[16'h3BE0] = 8'h00;
RAM[16'h3BE1] = 8'h00;
RAM[16'h3BE2] = 8'h00;
RAM[16'h3BE3] = 8'h00;
RAM[16'h3BE4] = 8'h00;
RAM[16'h3BE5] = 8'h00;
RAM[16'h3BE6] = 8'h00;
RAM[16'h3BE7] = 8'h00;
RAM[16'h3BE8] = 8'h00;
RAM[16'h3BE9] = 8'h00;
RAM[16'h3BEA] = 8'h00;
RAM[16'h3BEB] = 8'h00;
RAM[16'h3BEC] = 8'h00;
RAM[16'h3BED] = 8'h00;
RAM[16'h3BEE] = 8'h00;
RAM[16'h3BEF] = 8'h00;
RAM[16'h3BF0] = 8'h00;
RAM[16'h3BF1] = 8'h00;
RAM[16'h3BF2] = 8'h00;
RAM[16'h3BF3] = 8'h00;
RAM[16'h3BF4] = 8'h00;
RAM[16'h3BF5] = 8'h00;
RAM[16'h3BF6] = 8'h00;
RAM[16'h3BF7] = 8'h00;
RAM[16'h3BF8] = 8'h00;
RAM[16'h3BF9] = 8'h00;
RAM[16'h3BFA] = 8'h00;
RAM[16'h3BFB] = 8'h00;
RAM[16'h3BFC] = 8'h00;
RAM[16'h3BFD] = 8'h00;
RAM[16'h3BFE] = 8'h00;
RAM[16'h3BFF] = 8'h00;
RAM[16'h3C00] = 8'h00;
RAM[16'h3C01] = 8'h00;
RAM[16'h3C02] = 8'h00;
RAM[16'h3C03] = 8'h00;
RAM[16'h3C04] = 8'h00;
RAM[16'h3C05] = 8'h00;
RAM[16'h3C06] = 8'h00;
RAM[16'h3C07] = 8'h00;
RAM[16'h3C08] = 8'h00;
RAM[16'h3C09] = 8'h00;
RAM[16'h3C0A] = 8'h00;
RAM[16'h3C0B] = 8'h00;
RAM[16'h3C0C] = 8'h00;
RAM[16'h3C0D] = 8'h00;
RAM[16'h3C0E] = 8'h00;
RAM[16'h3C0F] = 8'h00;
RAM[16'h3C10] = 8'h00;
RAM[16'h3C11] = 8'h00;
RAM[16'h3C12] = 8'h00;
RAM[16'h3C13] = 8'h00;
RAM[16'h3C14] = 8'h00;
RAM[16'h3C15] = 8'h00;
RAM[16'h3C16] = 8'h00;
RAM[16'h3C17] = 8'h00;
RAM[16'h3C18] = 8'h00;
RAM[16'h3C19] = 8'h00;
RAM[16'h3C1A] = 8'h00;
RAM[16'h3C1B] = 8'h00;
RAM[16'h3C1C] = 8'h00;
RAM[16'h3C1D] = 8'h00;
RAM[16'h3C1E] = 8'h00;
RAM[16'h3C1F] = 8'h00;
RAM[16'h3C20] = 8'h00;
RAM[16'h3C21] = 8'h00;
RAM[16'h3C22] = 8'h00;
RAM[16'h3C23] = 8'h00;
RAM[16'h3C24] = 8'h00;
RAM[16'h3C25] = 8'h00;
RAM[16'h3C26] = 8'h00;
RAM[16'h3C27] = 8'h00;
RAM[16'h3C28] = 8'h00;
RAM[16'h3C29] = 8'h00;
RAM[16'h3C2A] = 8'h00;
RAM[16'h3C2B] = 8'h00;
RAM[16'h3C2C] = 8'h00;
RAM[16'h3C2D] = 8'h00;
RAM[16'h3C2E] = 8'h00;
RAM[16'h3C2F] = 8'h00;
RAM[16'h3C30] = 8'h00;
RAM[16'h3C31] = 8'h00;
RAM[16'h3C32] = 8'h00;
RAM[16'h3C33] = 8'h00;
RAM[16'h3C34] = 8'h00;
RAM[16'h3C35] = 8'h00;
RAM[16'h3C36] = 8'h00;
RAM[16'h3C37] = 8'h00;
RAM[16'h3C38] = 8'h00;
RAM[16'h3C39] = 8'h00;
RAM[16'h3C3A] = 8'h00;
RAM[16'h3C3B] = 8'h00;
RAM[16'h3C3C] = 8'h00;
RAM[16'h3C3D] = 8'h00;
RAM[16'h3C3E] = 8'h00;
RAM[16'h3C3F] = 8'h00;
RAM[16'h3C40] = 8'h00;
RAM[16'h3C41] = 8'h00;
RAM[16'h3C42] = 8'h00;
RAM[16'h3C43] = 8'h00;
RAM[16'h3C44] = 8'h00;
RAM[16'h3C45] = 8'h00;
RAM[16'h3C46] = 8'h00;
RAM[16'h3C47] = 8'h00;
RAM[16'h3C48] = 8'h00;
RAM[16'h3C49] = 8'h00;
RAM[16'h3C4A] = 8'h00;
RAM[16'h3C4B] = 8'h00;
RAM[16'h3C4C] = 8'h00;
RAM[16'h3C4D] = 8'h00;
RAM[16'h3C4E] = 8'h00;
RAM[16'h3C4F] = 8'h00;
RAM[16'h3C50] = 8'h00;
RAM[16'h3C51] = 8'h00;
RAM[16'h3C52] = 8'h00;
RAM[16'h3C53] = 8'h00;
RAM[16'h3C54] = 8'h00;
RAM[16'h3C55] = 8'h00;
RAM[16'h3C56] = 8'h00;
RAM[16'h3C57] = 8'h00;
RAM[16'h3C58] = 8'h00;
RAM[16'h3C59] = 8'h00;
RAM[16'h3C5A] = 8'h00;
RAM[16'h3C5B] = 8'h00;
RAM[16'h3C5C] = 8'h00;
RAM[16'h3C5D] = 8'h00;
RAM[16'h3C5E] = 8'h00;
RAM[16'h3C5F] = 8'h00;
RAM[16'h3C60] = 8'h00;
RAM[16'h3C61] = 8'h00;
RAM[16'h3C62] = 8'h00;
RAM[16'h3C63] = 8'h00;
RAM[16'h3C64] = 8'h00;
RAM[16'h3C65] = 8'h00;
RAM[16'h3C66] = 8'h00;
RAM[16'h3C67] = 8'h00;
RAM[16'h3C68] = 8'h00;
RAM[16'h3C69] = 8'h00;
RAM[16'h3C6A] = 8'h00;
RAM[16'h3C6B] = 8'h00;
RAM[16'h3C6C] = 8'h00;
RAM[16'h3C6D] = 8'h00;
RAM[16'h3C6E] = 8'h00;
RAM[16'h3C6F] = 8'h00;
RAM[16'h3C70] = 8'h00;
RAM[16'h3C71] = 8'h00;
RAM[16'h3C72] = 8'h00;
RAM[16'h3C73] = 8'h00;
RAM[16'h3C74] = 8'h00;
RAM[16'h3C75] = 8'h00;
RAM[16'h3C76] = 8'h00;
RAM[16'h3C77] = 8'h00;
RAM[16'h3C78] = 8'h00;
RAM[16'h3C79] = 8'h00;
RAM[16'h3C7A] = 8'h00;
RAM[16'h3C7B] = 8'h00;
RAM[16'h3C7C] = 8'h00;
RAM[16'h3C7D] = 8'h00;
RAM[16'h3C7E] = 8'h00;
RAM[16'h3C7F] = 8'h00;
RAM[16'h3C80] = 8'h00;
RAM[16'h3C81] = 8'h00;
RAM[16'h3C82] = 8'h00;
RAM[16'h3C83] = 8'h00;
RAM[16'h3C84] = 8'h00;
RAM[16'h3C85] = 8'h00;
RAM[16'h3C86] = 8'h00;
RAM[16'h3C87] = 8'h00;
RAM[16'h3C88] = 8'h00;
RAM[16'h3C89] = 8'h00;
RAM[16'h3C8A] = 8'h00;
RAM[16'h3C8B] = 8'h00;
RAM[16'h3C8C] = 8'h00;
RAM[16'h3C8D] = 8'h00;
RAM[16'h3C8E] = 8'h00;
RAM[16'h3C8F] = 8'h00;
RAM[16'h3C90] = 8'h00;
RAM[16'h3C91] = 8'h00;
RAM[16'h3C92] = 8'h00;
RAM[16'h3C93] = 8'h00;
RAM[16'h3C94] = 8'h00;
RAM[16'h3C95] = 8'h00;
RAM[16'h3C96] = 8'h00;
RAM[16'h3C97] = 8'h00;
RAM[16'h3C98] = 8'h00;
RAM[16'h3C99] = 8'h00;
RAM[16'h3C9A] = 8'h00;
RAM[16'h3C9B] = 8'h00;
RAM[16'h3C9C] = 8'h00;
RAM[16'h3C9D] = 8'h00;
RAM[16'h3C9E] = 8'h00;
RAM[16'h3C9F] = 8'h00;
RAM[16'h3CA0] = 8'h00;
RAM[16'h3CA1] = 8'h00;
RAM[16'h3CA2] = 8'h00;
RAM[16'h3CA3] = 8'h00;
RAM[16'h3CA4] = 8'h00;
RAM[16'h3CA5] = 8'h00;
RAM[16'h3CA6] = 8'h00;
RAM[16'h3CA7] = 8'h00;
RAM[16'h3CA8] = 8'h00;
RAM[16'h3CA9] = 8'h00;
RAM[16'h3CAA] = 8'h00;
RAM[16'h3CAB] = 8'h00;
RAM[16'h3CAC] = 8'h00;
RAM[16'h3CAD] = 8'h00;
RAM[16'h3CAE] = 8'h00;
RAM[16'h3CAF] = 8'h00;
RAM[16'h3CB0] = 8'h00;
RAM[16'h3CB1] = 8'h00;
RAM[16'h3CB2] = 8'h00;
RAM[16'h3CB3] = 8'h00;
RAM[16'h3CB4] = 8'h00;
RAM[16'h3CB5] = 8'h00;
RAM[16'h3CB6] = 8'h00;
RAM[16'h3CB7] = 8'h00;
RAM[16'h3CB8] = 8'h00;
RAM[16'h3CB9] = 8'h00;
RAM[16'h3CBA] = 8'h00;
RAM[16'h3CBB] = 8'h00;
RAM[16'h3CBC] = 8'h00;
RAM[16'h3CBD] = 8'h00;
RAM[16'h3CBE] = 8'h00;
RAM[16'h3CBF] = 8'h00;
RAM[16'h3CC0] = 8'h00;
RAM[16'h3CC1] = 8'h00;
RAM[16'h3CC2] = 8'h00;
RAM[16'h3CC3] = 8'h00;
RAM[16'h3CC4] = 8'h00;
RAM[16'h3CC5] = 8'h00;
RAM[16'h3CC6] = 8'h00;
RAM[16'h3CC7] = 8'h00;
RAM[16'h3CC8] = 8'h00;
RAM[16'h3CC9] = 8'h00;
RAM[16'h3CCA] = 8'h00;
RAM[16'h3CCB] = 8'h00;
RAM[16'h3CCC] = 8'h00;
RAM[16'h3CCD] = 8'h00;
RAM[16'h3CCE] = 8'h00;
RAM[16'h3CCF] = 8'h00;
RAM[16'h3CD0] = 8'h00;
RAM[16'h3CD1] = 8'h00;
RAM[16'h3CD2] = 8'h00;
RAM[16'h3CD3] = 8'h00;
RAM[16'h3CD4] = 8'h00;
RAM[16'h3CD5] = 8'h00;
RAM[16'h3CD6] = 8'h00;
RAM[16'h3CD7] = 8'h00;
RAM[16'h3CD8] = 8'h00;
RAM[16'h3CD9] = 8'h00;
RAM[16'h3CDA] = 8'h00;
RAM[16'h3CDB] = 8'h00;
RAM[16'h3CDC] = 8'h00;
RAM[16'h3CDD] = 8'h00;
RAM[16'h3CDE] = 8'h00;
RAM[16'h3CDF] = 8'h00;
RAM[16'h3CE0] = 8'h00;
RAM[16'h3CE1] = 8'h00;
RAM[16'h3CE2] = 8'h00;
RAM[16'h3CE3] = 8'h00;
RAM[16'h3CE4] = 8'h00;
RAM[16'h3CE5] = 8'h00;
RAM[16'h3CE6] = 8'h00;
RAM[16'h3CE7] = 8'h00;
RAM[16'h3CE8] = 8'h00;
RAM[16'h3CE9] = 8'h00;
RAM[16'h3CEA] = 8'h00;
RAM[16'h3CEB] = 8'h00;
RAM[16'h3CEC] = 8'h00;
RAM[16'h3CED] = 8'h00;
RAM[16'h3CEE] = 8'h00;
RAM[16'h3CEF] = 8'h00;
RAM[16'h3CF0] = 8'h00;
RAM[16'h3CF1] = 8'h00;
RAM[16'h3CF2] = 8'h00;
RAM[16'h3CF3] = 8'h00;
RAM[16'h3CF4] = 8'h00;
RAM[16'h3CF5] = 8'h00;
RAM[16'h3CF6] = 8'h00;
RAM[16'h3CF7] = 8'h00;
RAM[16'h3CF8] = 8'h00;
RAM[16'h3CF9] = 8'h00;
RAM[16'h3CFA] = 8'h00;
RAM[16'h3CFB] = 8'h00;
RAM[16'h3CFC] = 8'h00;
RAM[16'h3CFD] = 8'h00;
RAM[16'h3CFE] = 8'h00;
RAM[16'h3CFF] = 8'h00;
RAM[16'h3D00] = 8'h00;
RAM[16'h3D01] = 8'h00;
RAM[16'h3D02] = 8'h00;
RAM[16'h3D03] = 8'h00;
RAM[16'h3D04] = 8'h00;
RAM[16'h3D05] = 8'h00;
RAM[16'h3D06] = 8'h00;
RAM[16'h3D07] = 8'h00;
RAM[16'h3D08] = 8'h00;
RAM[16'h3D09] = 8'h00;
RAM[16'h3D0A] = 8'h00;
RAM[16'h3D0B] = 8'h00;
RAM[16'h3D0C] = 8'h00;
RAM[16'h3D0D] = 8'h00;
RAM[16'h3D0E] = 8'h00;
RAM[16'h3D0F] = 8'h00;
RAM[16'h3D10] = 8'h00;
RAM[16'h3D11] = 8'h00;
RAM[16'h3D12] = 8'h00;
RAM[16'h3D13] = 8'h00;
RAM[16'h3D14] = 8'h00;
RAM[16'h3D15] = 8'h00;
RAM[16'h3D16] = 8'h00;
RAM[16'h3D17] = 8'h00;
RAM[16'h3D18] = 8'h00;
RAM[16'h3D19] = 8'h00;
RAM[16'h3D1A] = 8'h00;
RAM[16'h3D1B] = 8'h00;
RAM[16'h3D1C] = 8'h00;
RAM[16'h3D1D] = 8'h00;
RAM[16'h3D1E] = 8'h00;
RAM[16'h3D1F] = 8'h00;
RAM[16'h3D20] = 8'h00;
RAM[16'h3D21] = 8'h00;
RAM[16'h3D22] = 8'h00;
RAM[16'h3D23] = 8'h00;
RAM[16'h3D24] = 8'h00;
RAM[16'h3D25] = 8'h00;
RAM[16'h3D26] = 8'h00;
RAM[16'h3D27] = 8'h00;
RAM[16'h3D28] = 8'h00;
RAM[16'h3D29] = 8'h00;
RAM[16'h3D2A] = 8'h00;
RAM[16'h3D2B] = 8'h00;
RAM[16'h3D2C] = 8'h00;
RAM[16'h3D2D] = 8'h00;
RAM[16'h3D2E] = 8'h00;
RAM[16'h3D2F] = 8'h00;
RAM[16'h3D30] = 8'h00;
RAM[16'h3D31] = 8'h00;
RAM[16'h3D32] = 8'h00;
RAM[16'h3D33] = 8'h00;
RAM[16'h3D34] = 8'h00;
RAM[16'h3D35] = 8'h00;
RAM[16'h3D36] = 8'h00;
RAM[16'h3D37] = 8'h00;
RAM[16'h3D38] = 8'h00;
RAM[16'h3D39] = 8'h00;
RAM[16'h3D3A] = 8'h00;
RAM[16'h3D3B] = 8'h00;
RAM[16'h3D3C] = 8'h00;
RAM[16'h3D3D] = 8'h00;
RAM[16'h3D3E] = 8'h00;
RAM[16'h3D3F] = 8'h00;
RAM[16'h3D40] = 8'h00;
RAM[16'h3D41] = 8'h00;
RAM[16'h3D42] = 8'h00;
RAM[16'h3D43] = 8'h00;
RAM[16'h3D44] = 8'h00;
RAM[16'h3D45] = 8'h00;
RAM[16'h3D46] = 8'h00;
RAM[16'h3D47] = 8'h00;
RAM[16'h3D48] = 8'h00;
RAM[16'h3D49] = 8'h00;
RAM[16'h3D4A] = 8'h00;
RAM[16'h3D4B] = 8'h00;
RAM[16'h3D4C] = 8'h00;
RAM[16'h3D4D] = 8'h00;
RAM[16'h3D4E] = 8'h00;
RAM[16'h3D4F] = 8'h00;
RAM[16'h3D50] = 8'h00;
RAM[16'h3D51] = 8'h00;
RAM[16'h3D52] = 8'h00;
RAM[16'h3D53] = 8'h00;
RAM[16'h3D54] = 8'h00;
RAM[16'h3D55] = 8'h00;
RAM[16'h3D56] = 8'h00;
RAM[16'h3D57] = 8'h00;
RAM[16'h3D58] = 8'h00;
RAM[16'h3D59] = 8'h00;
RAM[16'h3D5A] = 8'h00;
RAM[16'h3D5B] = 8'h00;
RAM[16'h3D5C] = 8'h00;
RAM[16'h3D5D] = 8'h00;
RAM[16'h3D5E] = 8'h00;
RAM[16'h3D5F] = 8'h00;
RAM[16'h3D60] = 8'h00;
RAM[16'h3D61] = 8'h00;
RAM[16'h3D62] = 8'h00;
RAM[16'h3D63] = 8'h00;
RAM[16'h3D64] = 8'h00;
RAM[16'h3D65] = 8'h00;
RAM[16'h3D66] = 8'h00;
RAM[16'h3D67] = 8'h00;
RAM[16'h3D68] = 8'h00;
RAM[16'h3D69] = 8'h00;
RAM[16'h3D6A] = 8'h00;
RAM[16'h3D6B] = 8'h00;
RAM[16'h3D6C] = 8'h00;
RAM[16'h3D6D] = 8'h00;
RAM[16'h3D6E] = 8'h00;
RAM[16'h3D6F] = 8'h00;
RAM[16'h3D70] = 8'h00;
RAM[16'h3D71] = 8'h00;
RAM[16'h3D72] = 8'h00;
RAM[16'h3D73] = 8'h00;
RAM[16'h3D74] = 8'h00;
RAM[16'h3D75] = 8'h00;
RAM[16'h3D76] = 8'h00;
RAM[16'h3D77] = 8'h00;
RAM[16'h3D78] = 8'h00;
RAM[16'h3D79] = 8'h00;
RAM[16'h3D7A] = 8'h00;
RAM[16'h3D7B] = 8'h00;
RAM[16'h3D7C] = 8'h00;
RAM[16'h3D7D] = 8'h00;
RAM[16'h3D7E] = 8'h00;
RAM[16'h3D7F] = 8'h00;
RAM[16'h3D80] = 8'h00;
RAM[16'h3D81] = 8'h00;
RAM[16'h3D82] = 8'h00;
RAM[16'h3D83] = 8'h00;
RAM[16'h3D84] = 8'h00;
RAM[16'h3D85] = 8'h00;
RAM[16'h3D86] = 8'h00;
RAM[16'h3D87] = 8'h00;
RAM[16'h3D88] = 8'h00;
RAM[16'h3D89] = 8'h00;
RAM[16'h3D8A] = 8'h00;
RAM[16'h3D8B] = 8'h00;
RAM[16'h3D8C] = 8'h00;
RAM[16'h3D8D] = 8'h00;
RAM[16'h3D8E] = 8'h00;
RAM[16'h3D8F] = 8'h00;
RAM[16'h3D90] = 8'h00;
RAM[16'h3D91] = 8'h00;
RAM[16'h3D92] = 8'h00;
RAM[16'h3D93] = 8'h00;
RAM[16'h3D94] = 8'h00;
RAM[16'h3D95] = 8'h00;
RAM[16'h3D96] = 8'h00;
RAM[16'h3D97] = 8'h00;
RAM[16'h3D98] = 8'h00;
RAM[16'h3D99] = 8'h00;
RAM[16'h3D9A] = 8'h00;
RAM[16'h3D9B] = 8'h00;
RAM[16'h3D9C] = 8'h00;
RAM[16'h3D9D] = 8'h00;
RAM[16'h3D9E] = 8'h00;
RAM[16'h3D9F] = 8'h00;
RAM[16'h3DA0] = 8'h00;
RAM[16'h3DA1] = 8'h00;
RAM[16'h3DA2] = 8'h00;
RAM[16'h3DA3] = 8'h00;
RAM[16'h3DA4] = 8'h00;
RAM[16'h3DA5] = 8'h00;
RAM[16'h3DA6] = 8'h00;
RAM[16'h3DA7] = 8'h00;
RAM[16'h3DA8] = 8'h00;
RAM[16'h3DA9] = 8'h00;
RAM[16'h3DAA] = 8'h00;
RAM[16'h3DAB] = 8'h00;
RAM[16'h3DAC] = 8'h00;
RAM[16'h3DAD] = 8'h00;
RAM[16'h3DAE] = 8'h00;
RAM[16'h3DAF] = 8'h00;
RAM[16'h3DB0] = 8'h00;
RAM[16'h3DB1] = 8'h00;
RAM[16'h3DB2] = 8'h00;
RAM[16'h3DB3] = 8'h00;
RAM[16'h3DB4] = 8'h00;
RAM[16'h3DB5] = 8'h00;
RAM[16'h3DB6] = 8'h00;
RAM[16'h3DB7] = 8'h00;
RAM[16'h3DB8] = 8'h00;
RAM[16'h3DB9] = 8'h00;
RAM[16'h3DBA] = 8'h00;
RAM[16'h3DBB] = 8'h00;
RAM[16'h3DBC] = 8'h00;
RAM[16'h3DBD] = 8'h00;
RAM[16'h3DBE] = 8'h00;
RAM[16'h3DBF] = 8'h00;
RAM[16'h3DC0] = 8'h00;
RAM[16'h3DC1] = 8'h00;
RAM[16'h3DC2] = 8'h00;
RAM[16'h3DC3] = 8'h00;
RAM[16'h3DC4] = 8'h00;
RAM[16'h3DC5] = 8'h00;
RAM[16'h3DC6] = 8'h00;
RAM[16'h3DC7] = 8'h00;
RAM[16'h3DC8] = 8'h00;
RAM[16'h3DC9] = 8'h00;
RAM[16'h3DCA] = 8'h00;
RAM[16'h3DCB] = 8'h00;
RAM[16'h3DCC] = 8'h00;
RAM[16'h3DCD] = 8'h00;
RAM[16'h3DCE] = 8'h00;
RAM[16'h3DCF] = 8'h00;
RAM[16'h3DD0] = 8'h00;
RAM[16'h3DD1] = 8'h00;
RAM[16'h3DD2] = 8'h00;
RAM[16'h3DD3] = 8'h00;
RAM[16'h3DD4] = 8'h00;
RAM[16'h3DD5] = 8'h00;
RAM[16'h3DD6] = 8'h00;
RAM[16'h3DD7] = 8'h00;
RAM[16'h3DD8] = 8'h00;
RAM[16'h3DD9] = 8'h00;
RAM[16'h3DDA] = 8'h00;
RAM[16'h3DDB] = 8'h00;
RAM[16'h3DDC] = 8'h00;
RAM[16'h3DDD] = 8'h00;
RAM[16'h3DDE] = 8'h00;
RAM[16'h3DDF] = 8'h00;
RAM[16'h3DE0] = 8'h00;
RAM[16'h3DE1] = 8'h00;
RAM[16'h3DE2] = 8'h00;
RAM[16'h3DE3] = 8'h00;
RAM[16'h3DE4] = 8'h00;
RAM[16'h3DE5] = 8'h00;
RAM[16'h3DE6] = 8'h00;
RAM[16'h3DE7] = 8'h00;
RAM[16'h3DE8] = 8'h00;
RAM[16'h3DE9] = 8'h00;
RAM[16'h3DEA] = 8'h00;
RAM[16'h3DEB] = 8'h00;
RAM[16'h3DEC] = 8'h00;
RAM[16'h3DED] = 8'h00;
RAM[16'h3DEE] = 8'h00;
RAM[16'h3DEF] = 8'h00;
RAM[16'h3DF0] = 8'h00;
RAM[16'h3DF1] = 8'h00;
RAM[16'h3DF2] = 8'h00;
RAM[16'h3DF3] = 8'h00;
RAM[16'h3DF4] = 8'h00;
RAM[16'h3DF5] = 8'h00;
RAM[16'h3DF6] = 8'h00;
RAM[16'h3DF7] = 8'h00;
RAM[16'h3DF8] = 8'h00;
RAM[16'h3DF9] = 8'h00;
RAM[16'h3DFA] = 8'h00;
RAM[16'h3DFB] = 8'h00;
RAM[16'h3DFC] = 8'h00;
RAM[16'h3DFD] = 8'h00;
RAM[16'h3DFE] = 8'h00;
RAM[16'h3DFF] = 8'h00;
RAM[16'h3E00] = 8'h00;
RAM[16'h3E01] = 8'h00;
RAM[16'h3E02] = 8'h00;
RAM[16'h3E03] = 8'h00;
RAM[16'h3E04] = 8'h00;
RAM[16'h3E05] = 8'h00;
RAM[16'h3E06] = 8'h00;
RAM[16'h3E07] = 8'h00;
RAM[16'h3E08] = 8'h00;
RAM[16'h3E09] = 8'h00;
RAM[16'h3E0A] = 8'h00;
RAM[16'h3E0B] = 8'h00;
RAM[16'h3E0C] = 8'h00;
RAM[16'h3E0D] = 8'h00;
RAM[16'h3E0E] = 8'h00;
RAM[16'h3E0F] = 8'h00;
RAM[16'h3E10] = 8'h00;
RAM[16'h3E11] = 8'h00;
RAM[16'h3E12] = 8'h00;
RAM[16'h3E13] = 8'h00;
RAM[16'h3E14] = 8'h00;
RAM[16'h3E15] = 8'h00;
RAM[16'h3E16] = 8'h00;
RAM[16'h3E17] = 8'h00;
RAM[16'h3E18] = 8'h00;
RAM[16'h3E19] = 8'h00;
RAM[16'h3E1A] = 8'h00;
RAM[16'h3E1B] = 8'h00;
RAM[16'h3E1C] = 8'h00;
RAM[16'h3E1D] = 8'h00;
RAM[16'h3E1E] = 8'h00;
RAM[16'h3E1F] = 8'h00;
RAM[16'h3E20] = 8'h00;
RAM[16'h3E21] = 8'h00;
RAM[16'h3E22] = 8'h00;
RAM[16'h3E23] = 8'h00;
RAM[16'h3E24] = 8'h00;
RAM[16'h3E25] = 8'h00;
RAM[16'h3E26] = 8'h00;
RAM[16'h3E27] = 8'h00;
RAM[16'h3E28] = 8'h00;
RAM[16'h3E29] = 8'h00;
RAM[16'h3E2A] = 8'h00;
RAM[16'h3E2B] = 8'h00;
RAM[16'h3E2C] = 8'h00;
RAM[16'h3E2D] = 8'h00;
RAM[16'h3E2E] = 8'h00;
RAM[16'h3E2F] = 8'h00;
RAM[16'h3E30] = 8'h00;
RAM[16'h3E31] = 8'h00;
RAM[16'h3E32] = 8'h00;
RAM[16'h3E33] = 8'h00;
RAM[16'h3E34] = 8'h00;
RAM[16'h3E35] = 8'h00;
RAM[16'h3E36] = 8'h00;
RAM[16'h3E37] = 8'h00;
RAM[16'h3E38] = 8'h00;
RAM[16'h3E39] = 8'h00;
RAM[16'h3E3A] = 8'h00;
RAM[16'h3E3B] = 8'h00;
RAM[16'h3E3C] = 8'h00;
RAM[16'h3E3D] = 8'h00;
RAM[16'h3E3E] = 8'h00;
RAM[16'h3E3F] = 8'h00;
RAM[16'h3E40] = 8'h00;
RAM[16'h3E41] = 8'h00;
RAM[16'h3E42] = 8'h00;
RAM[16'h3E43] = 8'h00;
RAM[16'h3E44] = 8'h00;
RAM[16'h3E45] = 8'h00;
RAM[16'h3E46] = 8'h00;
RAM[16'h3E47] = 8'h00;
RAM[16'h3E48] = 8'h00;
RAM[16'h3E49] = 8'h00;
RAM[16'h3E4A] = 8'h00;
RAM[16'h3E4B] = 8'h00;
RAM[16'h3E4C] = 8'h00;
RAM[16'h3E4D] = 8'h00;
RAM[16'h3E4E] = 8'h00;
RAM[16'h3E4F] = 8'h00;
RAM[16'h3E50] = 8'h00;
RAM[16'h3E51] = 8'h00;
RAM[16'h3E52] = 8'h00;
RAM[16'h3E53] = 8'h00;
RAM[16'h3E54] = 8'h00;
RAM[16'h3E55] = 8'h00;
RAM[16'h3E56] = 8'h00;
RAM[16'h3E57] = 8'h00;
RAM[16'h3E58] = 8'h00;
RAM[16'h3E59] = 8'h00;
RAM[16'h3E5A] = 8'h00;
RAM[16'h3E5B] = 8'h00;
RAM[16'h3E5C] = 8'h00;
RAM[16'h3E5D] = 8'h00;
RAM[16'h3E5E] = 8'h00;
RAM[16'h3E5F] = 8'h00;
RAM[16'h3E60] = 8'h00;
RAM[16'h3E61] = 8'h00;
RAM[16'h3E62] = 8'h00;
RAM[16'h3E63] = 8'h00;
RAM[16'h3E64] = 8'h00;
RAM[16'h3E65] = 8'h00;
RAM[16'h3E66] = 8'h00;
RAM[16'h3E67] = 8'h00;
RAM[16'h3E68] = 8'h00;
RAM[16'h3E69] = 8'h00;
RAM[16'h3E6A] = 8'h00;
RAM[16'h3E6B] = 8'h00;
RAM[16'h3E6C] = 8'h00;
RAM[16'h3E6D] = 8'h00;
RAM[16'h3E6E] = 8'h00;
RAM[16'h3E6F] = 8'h00;
RAM[16'h3E70] = 8'h00;
RAM[16'h3E71] = 8'h00;
RAM[16'h3E72] = 8'h00;
RAM[16'h3E73] = 8'h00;
RAM[16'h3E74] = 8'h00;
RAM[16'h3E75] = 8'h00;
RAM[16'h3E76] = 8'h00;
RAM[16'h3E77] = 8'h00;
RAM[16'h3E78] = 8'h00;
RAM[16'h3E79] = 8'h00;
RAM[16'h3E7A] = 8'h00;
RAM[16'h3E7B] = 8'h00;
RAM[16'h3E7C] = 8'h00;
RAM[16'h3E7D] = 8'h00;
RAM[16'h3E7E] = 8'h00;
RAM[16'h3E7F] = 8'h00;
RAM[16'h3E80] = 8'h00;
RAM[16'h3E81] = 8'h00;
RAM[16'h3E82] = 8'h00;
RAM[16'h3E83] = 8'h00;
RAM[16'h3E84] = 8'h00;
RAM[16'h3E85] = 8'h00;
RAM[16'h3E86] = 8'h00;
RAM[16'h3E87] = 8'h00;
RAM[16'h3E88] = 8'h00;
RAM[16'h3E89] = 8'h00;
RAM[16'h3E8A] = 8'h00;
RAM[16'h3E8B] = 8'h00;
RAM[16'h3E8C] = 8'h00;
RAM[16'h3E8D] = 8'h00;
RAM[16'h3E8E] = 8'h00;
RAM[16'h3E8F] = 8'h00;
RAM[16'h3E90] = 8'h00;
RAM[16'h3E91] = 8'h00;
RAM[16'h3E92] = 8'h00;
RAM[16'h3E93] = 8'h00;
RAM[16'h3E94] = 8'h00;
RAM[16'h3E95] = 8'h00;
RAM[16'h3E96] = 8'h00;
RAM[16'h3E97] = 8'h00;
RAM[16'h3E98] = 8'h00;
RAM[16'h3E99] = 8'h00;
RAM[16'h3E9A] = 8'h00;
RAM[16'h3E9B] = 8'h00;
RAM[16'h3E9C] = 8'h00;
RAM[16'h3E9D] = 8'h00;
RAM[16'h3E9E] = 8'h00;
RAM[16'h3E9F] = 8'h00;
RAM[16'h3EA0] = 8'h00;
RAM[16'h3EA1] = 8'h00;
RAM[16'h3EA2] = 8'h00;
RAM[16'h3EA3] = 8'h00;
RAM[16'h3EA4] = 8'h00;
RAM[16'h3EA5] = 8'h00;
RAM[16'h3EA6] = 8'h00;
RAM[16'h3EA7] = 8'h00;
RAM[16'h3EA8] = 8'h00;
RAM[16'h3EA9] = 8'h00;
RAM[16'h3EAA] = 8'h00;
RAM[16'h3EAB] = 8'h00;
RAM[16'h3EAC] = 8'h00;
RAM[16'h3EAD] = 8'h00;
RAM[16'h3EAE] = 8'h00;
RAM[16'h3EAF] = 8'h00;
RAM[16'h3EB0] = 8'h00;
RAM[16'h3EB1] = 8'h00;
RAM[16'h3EB2] = 8'h00;
RAM[16'h3EB3] = 8'h00;
RAM[16'h3EB4] = 8'h00;
RAM[16'h3EB5] = 8'h00;
RAM[16'h3EB6] = 8'h00;
RAM[16'h3EB7] = 8'h00;
RAM[16'h3EB8] = 8'h00;
RAM[16'h3EB9] = 8'h00;
RAM[16'h3EBA] = 8'h00;
RAM[16'h3EBB] = 8'h00;
RAM[16'h3EBC] = 8'h00;
RAM[16'h3EBD] = 8'h00;
RAM[16'h3EBE] = 8'h00;
RAM[16'h3EBF] = 8'h00;
RAM[16'h3EC0] = 8'h00;
RAM[16'h3EC1] = 8'h00;
RAM[16'h3EC2] = 8'h00;
RAM[16'h3EC3] = 8'h00;
RAM[16'h3EC4] = 8'h00;
RAM[16'h3EC5] = 8'h00;
RAM[16'h3EC6] = 8'h00;
RAM[16'h3EC7] = 8'h00;
RAM[16'h3EC8] = 8'h00;
RAM[16'h3EC9] = 8'h00;
RAM[16'h3ECA] = 8'h00;
RAM[16'h3ECB] = 8'h00;
RAM[16'h3ECC] = 8'h00;
RAM[16'h3ECD] = 8'h00;
RAM[16'h3ECE] = 8'h00;
RAM[16'h3ECF] = 8'h00;
RAM[16'h3ED0] = 8'h00;
RAM[16'h3ED1] = 8'h00;
RAM[16'h3ED2] = 8'h00;
RAM[16'h3ED3] = 8'h00;
RAM[16'h3ED4] = 8'h00;
RAM[16'h3ED5] = 8'h00;
RAM[16'h3ED6] = 8'h00;
RAM[16'h3ED7] = 8'h00;
RAM[16'h3ED8] = 8'h00;
RAM[16'h3ED9] = 8'h00;
RAM[16'h3EDA] = 8'h00;
RAM[16'h3EDB] = 8'h00;
RAM[16'h3EDC] = 8'h00;
RAM[16'h3EDD] = 8'h00;
RAM[16'h3EDE] = 8'h00;
RAM[16'h3EDF] = 8'h00;
RAM[16'h3EE0] = 8'h00;
RAM[16'h3EE1] = 8'h00;
RAM[16'h3EE2] = 8'h00;
RAM[16'h3EE3] = 8'h00;
RAM[16'h3EE4] = 8'h00;
RAM[16'h3EE5] = 8'h00;
RAM[16'h3EE6] = 8'h00;
RAM[16'h3EE7] = 8'h00;
RAM[16'h3EE8] = 8'h00;
RAM[16'h3EE9] = 8'h00;
RAM[16'h3EEA] = 8'h00;
RAM[16'h3EEB] = 8'h00;
RAM[16'h3EEC] = 8'h00;
RAM[16'h3EED] = 8'h00;
RAM[16'h3EEE] = 8'h00;
RAM[16'h3EEF] = 8'h00;
RAM[16'h3EF0] = 8'h00;
RAM[16'h3EF1] = 8'h00;
RAM[16'h3EF2] = 8'h00;
RAM[16'h3EF3] = 8'h00;
RAM[16'h3EF4] = 8'h00;
RAM[16'h3EF5] = 8'h00;
RAM[16'h3EF6] = 8'h00;
RAM[16'h3EF7] = 8'h00;
RAM[16'h3EF8] = 8'h00;
RAM[16'h3EF9] = 8'h00;
RAM[16'h3EFA] = 8'h00;
RAM[16'h3EFB] = 8'h00;
RAM[16'h3EFC] = 8'h00;
RAM[16'h3EFD] = 8'h00;
RAM[16'h3EFE] = 8'h00;
RAM[16'h3EFF] = 8'h00;
RAM[16'h3F00] = 8'h00;
RAM[16'h3F01] = 8'h00;
RAM[16'h3F02] = 8'h00;
RAM[16'h3F03] = 8'h00;
RAM[16'h3F04] = 8'h00;
RAM[16'h3F05] = 8'h00;
RAM[16'h3F06] = 8'h00;
RAM[16'h3F07] = 8'h00;
RAM[16'h3F08] = 8'h00;
RAM[16'h3F09] = 8'h00;
RAM[16'h3F0A] = 8'h00;
RAM[16'h3F0B] = 8'h00;
RAM[16'h3F0C] = 8'h00;
RAM[16'h3F0D] = 8'h00;
RAM[16'h3F0E] = 8'h00;
RAM[16'h3F0F] = 8'h00;
RAM[16'h3F10] = 8'h00;
RAM[16'h3F11] = 8'h00;
RAM[16'h3F12] = 8'h00;
RAM[16'h3F13] = 8'h00;
RAM[16'h3F14] = 8'h00;
RAM[16'h3F15] = 8'h00;
RAM[16'h3F16] = 8'h00;
RAM[16'h3F17] = 8'h00;
RAM[16'h3F18] = 8'h00;
RAM[16'h3F19] = 8'h00;
RAM[16'h3F1A] = 8'h00;
RAM[16'h3F1B] = 8'h00;
RAM[16'h3F1C] = 8'h00;
RAM[16'h3F1D] = 8'h00;
RAM[16'h3F1E] = 8'h00;
RAM[16'h3F1F] = 8'h00;
RAM[16'h3F20] = 8'h00;
RAM[16'h3F21] = 8'h00;
RAM[16'h3F22] = 8'h00;
RAM[16'h3F23] = 8'h00;
RAM[16'h3F24] = 8'h00;
RAM[16'h3F25] = 8'h00;
RAM[16'h3F26] = 8'h00;
RAM[16'h3F27] = 8'h00;
RAM[16'h3F28] = 8'h00;
RAM[16'h3F29] = 8'h00;
RAM[16'h3F2A] = 8'h00;
RAM[16'h3F2B] = 8'h00;
RAM[16'h3F2C] = 8'h00;
RAM[16'h3F2D] = 8'h00;
RAM[16'h3F2E] = 8'h00;
RAM[16'h3F2F] = 8'h00;
RAM[16'h3F30] = 8'h00;
RAM[16'h3F31] = 8'h00;
RAM[16'h3F32] = 8'h00;
RAM[16'h3F33] = 8'h00;
RAM[16'h3F34] = 8'h00;
RAM[16'h3F35] = 8'h00;
RAM[16'h3F36] = 8'h00;
RAM[16'h3F37] = 8'h00;
RAM[16'h3F38] = 8'h00;
RAM[16'h3F39] = 8'h00;
RAM[16'h3F3A] = 8'h00;
RAM[16'h3F3B] = 8'h00;
RAM[16'h3F3C] = 8'h00;
RAM[16'h3F3D] = 8'h00;
RAM[16'h3F3E] = 8'h00;
RAM[16'h3F3F] = 8'h00;
RAM[16'h3F40] = 8'h00;
RAM[16'h3F41] = 8'h00;
RAM[16'h3F42] = 8'h00;
RAM[16'h3F43] = 8'h00;
RAM[16'h3F44] = 8'h00;
RAM[16'h3F45] = 8'h00;
RAM[16'h3F46] = 8'h00;
RAM[16'h3F47] = 8'h00;
RAM[16'h3F48] = 8'h00;
RAM[16'h3F49] = 8'h00;
RAM[16'h3F4A] = 8'h00;
RAM[16'h3F4B] = 8'h00;
RAM[16'h3F4C] = 8'h00;
RAM[16'h3F4D] = 8'h00;
RAM[16'h3F4E] = 8'h00;
RAM[16'h3F4F] = 8'h00;
RAM[16'h3F50] = 8'h00;
RAM[16'h3F51] = 8'h00;
RAM[16'h3F52] = 8'h00;
RAM[16'h3F53] = 8'h00;
RAM[16'h3F54] = 8'h00;
RAM[16'h3F55] = 8'h00;
RAM[16'h3F56] = 8'h00;
RAM[16'h3F57] = 8'h00;
RAM[16'h3F58] = 8'h00;
RAM[16'h3F59] = 8'h00;
RAM[16'h3F5A] = 8'h00;
RAM[16'h3F5B] = 8'h00;
RAM[16'h3F5C] = 8'h00;
RAM[16'h3F5D] = 8'h00;
RAM[16'h3F5E] = 8'h00;
RAM[16'h3F5F] = 8'h00;
RAM[16'h3F60] = 8'h00;
RAM[16'h3F61] = 8'h00;
RAM[16'h3F62] = 8'h00;
RAM[16'h3F63] = 8'h00;
RAM[16'h3F64] = 8'h00;
RAM[16'h3F65] = 8'h00;
RAM[16'h3F66] = 8'h00;
RAM[16'h3F67] = 8'h00;
RAM[16'h3F68] = 8'h00;
RAM[16'h3F69] = 8'h00;
RAM[16'h3F6A] = 8'h00;
RAM[16'h3F6B] = 8'h00;
RAM[16'h3F6C] = 8'h00;
RAM[16'h3F6D] = 8'h00;
RAM[16'h3F6E] = 8'h00;
RAM[16'h3F6F] = 8'h00;
RAM[16'h3F70] = 8'h00;
RAM[16'h3F71] = 8'h00;
RAM[16'h3F72] = 8'h00;
RAM[16'h3F73] = 8'h00;
RAM[16'h3F74] = 8'h00;
RAM[16'h3F75] = 8'h00;
RAM[16'h3F76] = 8'h00;
RAM[16'h3F77] = 8'h00;
RAM[16'h3F78] = 8'h00;
RAM[16'h3F79] = 8'h00;
RAM[16'h3F7A] = 8'h00;
RAM[16'h3F7B] = 8'h00;
RAM[16'h3F7C] = 8'h00;
RAM[16'h3F7D] = 8'h00;
RAM[16'h3F7E] = 8'h00;
RAM[16'h3F7F] = 8'h00;
RAM[16'h3F80] = 8'h00;
RAM[16'h3F81] = 8'h00;
RAM[16'h3F82] = 8'h00;
RAM[16'h3F83] = 8'h00;
RAM[16'h3F84] = 8'h00;
RAM[16'h3F85] = 8'h00;
RAM[16'h3F86] = 8'h00;
RAM[16'h3F87] = 8'h00;
RAM[16'h3F88] = 8'h00;
RAM[16'h3F89] = 8'h00;
RAM[16'h3F8A] = 8'h00;
RAM[16'h3F8B] = 8'h00;
RAM[16'h3F8C] = 8'h00;
RAM[16'h3F8D] = 8'h00;
RAM[16'h3F8E] = 8'h00;
RAM[16'h3F8F] = 8'h00;
RAM[16'h3F90] = 8'h00;
RAM[16'h3F91] = 8'h00;
RAM[16'h3F92] = 8'h00;
RAM[16'h3F93] = 8'h00;
RAM[16'h3F94] = 8'h00;
RAM[16'h3F95] = 8'h00;
RAM[16'h3F96] = 8'h00;
RAM[16'h3F97] = 8'h00;
RAM[16'h3F98] = 8'h00;
RAM[16'h3F99] = 8'h00;
RAM[16'h3F9A] = 8'h00;
RAM[16'h3F9B] = 8'h00;
RAM[16'h3F9C] = 8'h00;
RAM[16'h3F9D] = 8'h00;
RAM[16'h3F9E] = 8'h00;
RAM[16'h3F9F] = 8'h00;
RAM[16'h3FA0] = 8'h00;
RAM[16'h3FA1] = 8'h00;
RAM[16'h3FA2] = 8'h00;
RAM[16'h3FA3] = 8'h00;
RAM[16'h3FA4] = 8'h00;
RAM[16'h3FA5] = 8'h00;
RAM[16'h3FA6] = 8'h00;
RAM[16'h3FA7] = 8'h00;
RAM[16'h3FA8] = 8'h00;
RAM[16'h3FA9] = 8'h00;
RAM[16'h3FAA] = 8'h00;
RAM[16'h3FAB] = 8'h00;
RAM[16'h3FAC] = 8'h00;
RAM[16'h3FAD] = 8'h00;
RAM[16'h3FAE] = 8'h00;
RAM[16'h3FAF] = 8'h00;
RAM[16'h3FB0] = 8'h00;
RAM[16'h3FB1] = 8'h00;
RAM[16'h3FB2] = 8'h00;
RAM[16'h3FB3] = 8'h00;
RAM[16'h3FB4] = 8'h00;
RAM[16'h3FB5] = 8'h00;
RAM[16'h3FB6] = 8'h00;
RAM[16'h3FB7] = 8'h00;
RAM[16'h3FB8] = 8'h00;
RAM[16'h3FB9] = 8'h00;
RAM[16'h3FBA] = 8'h00;
RAM[16'h3FBB] = 8'h00;
RAM[16'h3FBC] = 8'h00;
RAM[16'h3FBD] = 8'h00;
RAM[16'h3FBE] = 8'h00;
RAM[16'h3FBF] = 8'h00;
RAM[16'h3FC0] = 8'h00;
RAM[16'h3FC1] = 8'h00;
RAM[16'h3FC2] = 8'h00;
RAM[16'h3FC3] = 8'h00;
RAM[16'h3FC4] = 8'h00;
RAM[16'h3FC5] = 8'h00;
RAM[16'h3FC6] = 8'h00;
RAM[16'h3FC7] = 8'h00;
RAM[16'h3FC8] = 8'h00;
RAM[16'h3FC9] = 8'h00;
RAM[16'h3FCA] = 8'h00;
RAM[16'h3FCB] = 8'h00;
RAM[16'h3FCC] = 8'h00;
RAM[16'h3FCD] = 8'h00;
RAM[16'h3FCE] = 8'h00;
RAM[16'h3FCF] = 8'h00;
RAM[16'h3FD0] = 8'h00;
RAM[16'h3FD1] = 8'h00;
RAM[16'h3FD2] = 8'h00;
RAM[16'h3FD3] = 8'h00;
RAM[16'h3FD4] = 8'h00;
RAM[16'h3FD5] = 8'h00;
RAM[16'h3FD6] = 8'h00;
RAM[16'h3FD7] = 8'h00;
RAM[16'h3FD8] = 8'h00;
RAM[16'h3FD9] = 8'h00;
RAM[16'h3FDA] = 8'h00;
RAM[16'h3FDB] = 8'h00;
RAM[16'h3FDC] = 8'h00;
RAM[16'h3FDD] = 8'h00;
RAM[16'h3FDE] = 8'h00;
RAM[16'h3FDF] = 8'h00;
RAM[16'h3FE0] = 8'h00;
RAM[16'h3FE1] = 8'h00;
RAM[16'h3FE2] = 8'h00;
RAM[16'h3FE3] = 8'h00;
RAM[16'h3FE4] = 8'h00;
RAM[16'h3FE5] = 8'h00;
RAM[16'h3FE6] = 8'h00;
RAM[16'h3FE7] = 8'h00;
RAM[16'h3FE8] = 8'h00;
RAM[16'h3FE9] = 8'h00;
RAM[16'h3FEA] = 8'h00;
RAM[16'h3FEB] = 8'h00;
RAM[16'h3FEC] = 8'h00;
RAM[16'h3FED] = 8'h00;
RAM[16'h3FEE] = 8'h00;
RAM[16'h3FEF] = 8'h00;
RAM[16'h3FF0] = 8'h00;
RAM[16'h3FF1] = 8'h00;
RAM[16'h3FF2] = 8'h00;
RAM[16'h3FF3] = 8'h00;
RAM[16'h3FF4] = 8'h00;
RAM[16'h3FF5] = 8'h00;
RAM[16'h3FF6] = 8'h00;
RAM[16'h3FF7] = 8'h00;
RAM[16'h3FF8] = 8'h00;
RAM[16'h3FF9] = 8'h00;
RAM[16'h3FFA] = 8'h00;
RAM[16'h3FFB] = 8'h00;
RAM[16'h3FFC] = 8'h00;
RAM[16'h3FFD] = 8'h00;
RAM[16'h3FFE] = 8'h00;
RAM[16'h3FFF] = 8'h00;
RAM[16'h4000] = 8'h00;
RAM[16'h4001] = 8'h00;
RAM[16'h4002] = 8'h00;
RAM[16'h4003] = 8'h00;
RAM[16'h4004] = 8'h00;
RAM[16'h4005] = 8'h00;
RAM[16'h4006] = 8'h00;
RAM[16'h4007] = 8'h00;
RAM[16'h4008] = 8'h00;
RAM[16'h4009] = 8'h00;
RAM[16'h400A] = 8'h00;
RAM[16'h400B] = 8'h00;
RAM[16'h400C] = 8'h00;
RAM[16'h400D] = 8'h00;
RAM[16'h400E] = 8'h00;
RAM[16'h400F] = 8'h00;
RAM[16'h4010] = 8'h00;
RAM[16'h4011] = 8'h00;
RAM[16'h4012] = 8'h00;
RAM[16'h4013] = 8'h00;
RAM[16'h4014] = 8'h00;
RAM[16'h4015] = 8'h00;
RAM[16'h4016] = 8'h00;
RAM[16'h4017] = 8'h00;
RAM[16'h4018] = 8'h00;
RAM[16'h4019] = 8'h00;
RAM[16'h401A] = 8'h00;
RAM[16'h401B] = 8'h00;
RAM[16'h401C] = 8'h00;
RAM[16'h401D] = 8'h00;
RAM[16'h401E] = 8'h00;
RAM[16'h401F] = 8'h00;
RAM[16'h4020] = 8'h00;
RAM[16'h4021] = 8'h00;
RAM[16'h4022] = 8'h00;
RAM[16'h4023] = 8'h00;
RAM[16'h4024] = 8'h00;
RAM[16'h4025] = 8'h00;
RAM[16'h4026] = 8'h00;
RAM[16'h4027] = 8'h00;
RAM[16'h4028] = 8'h00;
RAM[16'h4029] = 8'h00;
RAM[16'h402A] = 8'h00;
RAM[16'h402B] = 8'h00;
RAM[16'h402C] = 8'h00;
RAM[16'h402D] = 8'h00;
RAM[16'h402E] = 8'h00;
RAM[16'h402F] = 8'h00;
RAM[16'h4030] = 8'h00;
RAM[16'h4031] = 8'h00;
RAM[16'h4032] = 8'h00;
RAM[16'h4033] = 8'h00;
RAM[16'h4034] = 8'h00;
RAM[16'h4035] = 8'h00;
RAM[16'h4036] = 8'h00;
RAM[16'h4037] = 8'h00;
RAM[16'h4038] = 8'h00;
RAM[16'h4039] = 8'h00;
RAM[16'h403A] = 8'h00;
RAM[16'h403B] = 8'h00;
RAM[16'h403C] = 8'h00;
RAM[16'h403D] = 8'h00;
RAM[16'h403E] = 8'h00;
RAM[16'h403F] = 8'h00;
RAM[16'h4040] = 8'h00;
RAM[16'h4041] = 8'h00;
RAM[16'h4042] = 8'h00;
RAM[16'h4043] = 8'h00;
RAM[16'h4044] = 8'h00;
RAM[16'h4045] = 8'h00;
RAM[16'h4046] = 8'h00;
RAM[16'h4047] = 8'h00;
RAM[16'h4048] = 8'h00;
RAM[16'h4049] = 8'h00;
RAM[16'h404A] = 8'h00;
RAM[16'h404B] = 8'h00;
RAM[16'h404C] = 8'h00;
RAM[16'h404D] = 8'h00;
RAM[16'h404E] = 8'h00;
RAM[16'h404F] = 8'h00;
RAM[16'h4050] = 8'h00;
RAM[16'h4051] = 8'h00;
RAM[16'h4052] = 8'h00;
RAM[16'h4053] = 8'h00;
RAM[16'h4054] = 8'h00;
RAM[16'h4055] = 8'h00;
RAM[16'h4056] = 8'h00;
RAM[16'h4057] = 8'h00;
RAM[16'h4058] = 8'h00;
RAM[16'h4059] = 8'h00;
RAM[16'h405A] = 8'h00;
RAM[16'h405B] = 8'h00;
RAM[16'h405C] = 8'h00;
RAM[16'h405D] = 8'h00;
RAM[16'h405E] = 8'h00;
RAM[16'h405F] = 8'h00;
RAM[16'h4060] = 8'h00;
RAM[16'h4061] = 8'h00;
RAM[16'h4062] = 8'h00;
RAM[16'h4063] = 8'h00;
RAM[16'h4064] = 8'h00;
RAM[16'h4065] = 8'h00;
RAM[16'h4066] = 8'h00;
RAM[16'h4067] = 8'h00;
RAM[16'h4068] = 8'h00;
RAM[16'h4069] = 8'h00;
RAM[16'h406A] = 8'h00;
RAM[16'h406B] = 8'h00;
RAM[16'h406C] = 8'h00;
RAM[16'h406D] = 8'h00;
RAM[16'h406E] = 8'h00;
RAM[16'h406F] = 8'h00;
RAM[16'h4070] = 8'h00;
RAM[16'h4071] = 8'h00;
RAM[16'h4072] = 8'h00;
RAM[16'h4073] = 8'h00;
RAM[16'h4074] = 8'h00;
RAM[16'h4075] = 8'h00;
RAM[16'h4076] = 8'h00;
RAM[16'h4077] = 8'h00;
RAM[16'h4078] = 8'h00;
RAM[16'h4079] = 8'h00;
RAM[16'h407A] = 8'h00;
RAM[16'h407B] = 8'h00;
RAM[16'h407C] = 8'h00;
RAM[16'h407D] = 8'h00;
RAM[16'h407E] = 8'h00;
RAM[16'h407F] = 8'h00;
RAM[16'h4080] = 8'h00;
RAM[16'h4081] = 8'h00;
RAM[16'h4082] = 8'h00;
RAM[16'h4083] = 8'h00;
RAM[16'h4084] = 8'h00;
RAM[16'h4085] = 8'h00;
RAM[16'h4086] = 8'h00;
RAM[16'h4087] = 8'h00;
RAM[16'h4088] = 8'h00;
RAM[16'h4089] = 8'h00;
RAM[16'h408A] = 8'h00;
RAM[16'h408B] = 8'h00;
RAM[16'h408C] = 8'h00;
RAM[16'h408D] = 8'h00;
RAM[16'h408E] = 8'h00;
RAM[16'h408F] = 8'h00;
RAM[16'h4090] = 8'h00;
RAM[16'h4091] = 8'h00;
RAM[16'h4092] = 8'h00;
RAM[16'h4093] = 8'h00;
RAM[16'h4094] = 8'h00;
RAM[16'h4095] = 8'h00;
RAM[16'h4096] = 8'h00;
RAM[16'h4097] = 8'h00;
RAM[16'h4098] = 8'h00;
RAM[16'h4099] = 8'h00;
RAM[16'h409A] = 8'h00;
RAM[16'h409B] = 8'h00;
RAM[16'h409C] = 8'h00;
RAM[16'h409D] = 8'h00;
RAM[16'h409E] = 8'h00;
RAM[16'h409F] = 8'h00;
RAM[16'h40A0] = 8'h00;
RAM[16'h40A1] = 8'h00;
RAM[16'h40A2] = 8'h00;
RAM[16'h40A3] = 8'h00;
RAM[16'h40A4] = 8'h00;
RAM[16'h40A5] = 8'h00;
RAM[16'h40A6] = 8'h00;
RAM[16'h40A7] = 8'h00;
RAM[16'h40A8] = 8'h00;
RAM[16'h40A9] = 8'h00;
RAM[16'h40AA] = 8'h00;
RAM[16'h40AB] = 8'h00;
RAM[16'h40AC] = 8'h00;
RAM[16'h40AD] = 8'h00;
RAM[16'h40AE] = 8'h00;
RAM[16'h40AF] = 8'h00;
RAM[16'h40B0] = 8'h00;
RAM[16'h40B1] = 8'h00;
RAM[16'h40B2] = 8'h00;
RAM[16'h40B3] = 8'h00;
RAM[16'h40B4] = 8'h00;
RAM[16'h40B5] = 8'h00;
RAM[16'h40B6] = 8'h00;
RAM[16'h40B7] = 8'h00;
RAM[16'h40B8] = 8'h00;
RAM[16'h40B9] = 8'h00;
RAM[16'h40BA] = 8'h00;
RAM[16'h40BB] = 8'h00;
RAM[16'h40BC] = 8'h00;
RAM[16'h40BD] = 8'h00;
RAM[16'h40BE] = 8'h00;
RAM[16'h40BF] = 8'h00;
RAM[16'h40C0] = 8'h00;
RAM[16'h40C1] = 8'h00;
RAM[16'h40C2] = 8'h00;
RAM[16'h40C3] = 8'h00;
RAM[16'h40C4] = 8'h00;
RAM[16'h40C5] = 8'h00;
RAM[16'h40C6] = 8'h00;
RAM[16'h40C7] = 8'h00;
RAM[16'h40C8] = 8'h00;
RAM[16'h40C9] = 8'h00;
RAM[16'h40CA] = 8'h00;
RAM[16'h40CB] = 8'h00;
RAM[16'h40CC] = 8'h00;
RAM[16'h40CD] = 8'h00;
RAM[16'h40CE] = 8'h00;
RAM[16'h40CF] = 8'h00;
RAM[16'h40D0] = 8'h00;
RAM[16'h40D1] = 8'h00;
RAM[16'h40D2] = 8'h00;
RAM[16'h40D3] = 8'h00;
RAM[16'h40D4] = 8'h00;
RAM[16'h40D5] = 8'h00;
RAM[16'h40D6] = 8'h00;
RAM[16'h40D7] = 8'h00;
RAM[16'h40D8] = 8'h00;
RAM[16'h40D9] = 8'h00;
RAM[16'h40DA] = 8'h00;
RAM[16'h40DB] = 8'h00;
RAM[16'h40DC] = 8'h00;
RAM[16'h40DD] = 8'h00;
RAM[16'h40DE] = 8'h00;
RAM[16'h40DF] = 8'h00;
RAM[16'h40E0] = 8'h00;
RAM[16'h40E1] = 8'h00;
RAM[16'h40E2] = 8'h00;
RAM[16'h40E3] = 8'h00;
RAM[16'h40E4] = 8'h00;
RAM[16'h40E5] = 8'h00;
RAM[16'h40E6] = 8'h00;
RAM[16'h40E7] = 8'h00;
RAM[16'h40E8] = 8'h00;
RAM[16'h40E9] = 8'h00;
RAM[16'h40EA] = 8'h00;
RAM[16'h40EB] = 8'h00;
RAM[16'h40EC] = 8'h00;
RAM[16'h40ED] = 8'h00;
RAM[16'h40EE] = 8'h00;
RAM[16'h40EF] = 8'h00;
RAM[16'h40F0] = 8'h00;
RAM[16'h40F1] = 8'h00;
RAM[16'h40F2] = 8'h00;
RAM[16'h40F3] = 8'h00;
RAM[16'h40F4] = 8'h00;
RAM[16'h40F5] = 8'h00;
RAM[16'h40F6] = 8'h00;
RAM[16'h40F7] = 8'h00;
RAM[16'h40F8] = 8'h00;
RAM[16'h40F9] = 8'h00;
RAM[16'h40FA] = 8'h00;
RAM[16'h40FB] = 8'h00;
RAM[16'h40FC] = 8'h00;
RAM[16'h40FD] = 8'h00;
RAM[16'h40FE] = 8'h00;
RAM[16'h40FF] = 8'h00;
RAM[16'h4100] = 8'h00;
RAM[16'h4101] = 8'h00;
RAM[16'h4102] = 8'h00;
RAM[16'h4103] = 8'h00;
RAM[16'h4104] = 8'h00;
RAM[16'h4105] = 8'h00;
RAM[16'h4106] = 8'h00;
RAM[16'h4107] = 8'h00;
RAM[16'h4108] = 8'h00;
RAM[16'h4109] = 8'h00;
RAM[16'h410A] = 8'h00;
RAM[16'h410B] = 8'h00;
RAM[16'h410C] = 8'h00;
RAM[16'h410D] = 8'h00;
RAM[16'h410E] = 8'h00;
RAM[16'h410F] = 8'h00;
RAM[16'h4110] = 8'h00;
RAM[16'h4111] = 8'h00;
RAM[16'h4112] = 8'h00;
RAM[16'h4113] = 8'h00;
RAM[16'h4114] = 8'h00;
RAM[16'h4115] = 8'h00;
RAM[16'h4116] = 8'h00;
RAM[16'h4117] = 8'h00;
RAM[16'h4118] = 8'h00;
RAM[16'h4119] = 8'h00;
RAM[16'h411A] = 8'h00;
RAM[16'h411B] = 8'h00;
RAM[16'h411C] = 8'h00;
RAM[16'h411D] = 8'h00;
RAM[16'h411E] = 8'h00;
RAM[16'h411F] = 8'h00;
RAM[16'h4120] = 8'h00;
RAM[16'h4121] = 8'h00;
RAM[16'h4122] = 8'h00;
RAM[16'h4123] = 8'h00;
RAM[16'h4124] = 8'h00;
RAM[16'h4125] = 8'h00;
RAM[16'h4126] = 8'h00;
RAM[16'h4127] = 8'h00;
RAM[16'h4128] = 8'h00;
RAM[16'h4129] = 8'h00;
RAM[16'h412A] = 8'h00;
RAM[16'h412B] = 8'h00;
RAM[16'h412C] = 8'h00;
RAM[16'h412D] = 8'h00;
RAM[16'h412E] = 8'h00;
RAM[16'h412F] = 8'h00;
RAM[16'h4130] = 8'h00;
RAM[16'h4131] = 8'h00;
RAM[16'h4132] = 8'h00;
RAM[16'h4133] = 8'h00;
RAM[16'h4134] = 8'h00;
RAM[16'h4135] = 8'h00;
RAM[16'h4136] = 8'h00;
RAM[16'h4137] = 8'h00;
RAM[16'h4138] = 8'h00;
RAM[16'h4139] = 8'h00;
RAM[16'h413A] = 8'h00;
RAM[16'h413B] = 8'h00;
RAM[16'h413C] = 8'h00;
RAM[16'h413D] = 8'h00;
RAM[16'h413E] = 8'h00;
RAM[16'h413F] = 8'h00;
RAM[16'h4140] = 8'h00;
RAM[16'h4141] = 8'h00;
RAM[16'h4142] = 8'h00;
RAM[16'h4143] = 8'h00;
RAM[16'h4144] = 8'h00;
RAM[16'h4145] = 8'h00;
RAM[16'h4146] = 8'h00;
RAM[16'h4147] = 8'h00;
RAM[16'h4148] = 8'h00;
RAM[16'h4149] = 8'h00;
RAM[16'h414A] = 8'h00;
RAM[16'h414B] = 8'h00;
RAM[16'h414C] = 8'h00;
RAM[16'h414D] = 8'h00;
RAM[16'h414E] = 8'h00;
RAM[16'h414F] = 8'h00;
RAM[16'h4150] = 8'h00;
RAM[16'h4151] = 8'h00;
RAM[16'h4152] = 8'h00;
RAM[16'h4153] = 8'h00;
RAM[16'h4154] = 8'h00;
RAM[16'h4155] = 8'h00;
RAM[16'h4156] = 8'h00;
RAM[16'h4157] = 8'h00;
RAM[16'h4158] = 8'h00;
RAM[16'h4159] = 8'h00;
RAM[16'h415A] = 8'h00;
RAM[16'h415B] = 8'h00;
RAM[16'h415C] = 8'h00;
RAM[16'h415D] = 8'h00;
RAM[16'h415E] = 8'h00;
RAM[16'h415F] = 8'h00;
RAM[16'h4160] = 8'h00;
RAM[16'h4161] = 8'h00;
RAM[16'h4162] = 8'h00;
RAM[16'h4163] = 8'h00;
RAM[16'h4164] = 8'h00;
RAM[16'h4165] = 8'h00;
RAM[16'h4166] = 8'h00;
RAM[16'h4167] = 8'h00;
RAM[16'h4168] = 8'h00;
RAM[16'h4169] = 8'h00;
RAM[16'h416A] = 8'h00;
RAM[16'h416B] = 8'h00;
RAM[16'h416C] = 8'h00;
RAM[16'h416D] = 8'h00;
RAM[16'h416E] = 8'h00;
RAM[16'h416F] = 8'h00;
RAM[16'h4170] = 8'h00;
RAM[16'h4171] = 8'h00;
RAM[16'h4172] = 8'h00;
RAM[16'h4173] = 8'h00;
RAM[16'h4174] = 8'h00;
RAM[16'h4175] = 8'h00;
RAM[16'h4176] = 8'h00;
RAM[16'h4177] = 8'h00;
RAM[16'h4178] = 8'h00;
RAM[16'h4179] = 8'h00;
RAM[16'h417A] = 8'h00;
RAM[16'h417B] = 8'h00;
RAM[16'h417C] = 8'h00;
RAM[16'h417D] = 8'h00;
RAM[16'h417E] = 8'h00;
RAM[16'h417F] = 8'h00;
RAM[16'h4180] = 8'h00;
RAM[16'h4181] = 8'h00;
RAM[16'h4182] = 8'h00;
RAM[16'h4183] = 8'h00;
RAM[16'h4184] = 8'h00;
RAM[16'h4185] = 8'h00;
RAM[16'h4186] = 8'h00;
RAM[16'h4187] = 8'h00;
RAM[16'h4188] = 8'h00;
RAM[16'h4189] = 8'h00;
RAM[16'h418A] = 8'h00;
RAM[16'h418B] = 8'h00;
RAM[16'h418C] = 8'h00;
RAM[16'h418D] = 8'h00;
RAM[16'h418E] = 8'h00;
RAM[16'h418F] = 8'h00;
RAM[16'h4190] = 8'h00;
RAM[16'h4191] = 8'h00;
RAM[16'h4192] = 8'h00;
RAM[16'h4193] = 8'h00;
RAM[16'h4194] = 8'h00;
RAM[16'h4195] = 8'h00;
RAM[16'h4196] = 8'h00;
RAM[16'h4197] = 8'h00;
RAM[16'h4198] = 8'h00;
RAM[16'h4199] = 8'h00;
RAM[16'h419A] = 8'h00;
RAM[16'h419B] = 8'h00;
RAM[16'h419C] = 8'h00;
RAM[16'h419D] = 8'h00;
RAM[16'h419E] = 8'h00;
RAM[16'h419F] = 8'h00;
RAM[16'h41A0] = 8'h00;
RAM[16'h41A1] = 8'h00;
RAM[16'h41A2] = 8'h00;
RAM[16'h41A3] = 8'h00;
RAM[16'h41A4] = 8'h00;
RAM[16'h41A5] = 8'h00;
RAM[16'h41A6] = 8'h00;
RAM[16'h41A7] = 8'h00;
RAM[16'h41A8] = 8'h00;
RAM[16'h41A9] = 8'h00;
RAM[16'h41AA] = 8'h00;
RAM[16'h41AB] = 8'h00;
RAM[16'h41AC] = 8'h00;
RAM[16'h41AD] = 8'h00;
RAM[16'h41AE] = 8'h00;
RAM[16'h41AF] = 8'h00;
RAM[16'h41B0] = 8'h00;
RAM[16'h41B1] = 8'h00;
RAM[16'h41B2] = 8'h00;
RAM[16'h41B3] = 8'h00;
RAM[16'h41B4] = 8'h00;
RAM[16'h41B5] = 8'h00;
RAM[16'h41B6] = 8'h00;
RAM[16'h41B7] = 8'h00;
RAM[16'h41B8] = 8'h00;
RAM[16'h41B9] = 8'h00;
RAM[16'h41BA] = 8'h00;
RAM[16'h41BB] = 8'h00;
RAM[16'h41BC] = 8'h00;
RAM[16'h41BD] = 8'h00;
RAM[16'h41BE] = 8'h00;
RAM[16'h41BF] = 8'h00;
RAM[16'h41C0] = 8'h00;
RAM[16'h41C1] = 8'h00;
RAM[16'h41C2] = 8'h00;
RAM[16'h41C3] = 8'h00;
RAM[16'h41C4] = 8'h00;
RAM[16'h41C5] = 8'h00;
RAM[16'h41C6] = 8'h00;
RAM[16'h41C7] = 8'h00;
RAM[16'h41C8] = 8'h00;
RAM[16'h41C9] = 8'h00;
RAM[16'h41CA] = 8'h00;
RAM[16'h41CB] = 8'h00;
RAM[16'h41CC] = 8'h00;
RAM[16'h41CD] = 8'h00;
RAM[16'h41CE] = 8'h00;
RAM[16'h41CF] = 8'h00;
RAM[16'h41D0] = 8'h00;
RAM[16'h41D1] = 8'h00;
RAM[16'h41D2] = 8'h00;
RAM[16'h41D3] = 8'h00;
RAM[16'h41D4] = 8'h00;
RAM[16'h41D5] = 8'h00;
RAM[16'h41D6] = 8'h00;
RAM[16'h41D7] = 8'h00;
RAM[16'h41D8] = 8'h00;
RAM[16'h41D9] = 8'h00;
RAM[16'h41DA] = 8'h00;
RAM[16'h41DB] = 8'h00;
RAM[16'h41DC] = 8'h00;
RAM[16'h41DD] = 8'h00;
RAM[16'h41DE] = 8'h00;
RAM[16'h41DF] = 8'h00;
RAM[16'h41E0] = 8'h00;
RAM[16'h41E1] = 8'h00;
RAM[16'h41E2] = 8'h00;
RAM[16'h41E3] = 8'h00;
RAM[16'h41E4] = 8'h00;
RAM[16'h41E5] = 8'h00;
RAM[16'h41E6] = 8'h00;
RAM[16'h41E7] = 8'h00;
RAM[16'h41E8] = 8'h00;
RAM[16'h41E9] = 8'h00;
RAM[16'h41EA] = 8'h00;
RAM[16'h41EB] = 8'h00;
RAM[16'h41EC] = 8'h00;
RAM[16'h41ED] = 8'h00;
RAM[16'h41EE] = 8'h00;
RAM[16'h41EF] = 8'h00;
RAM[16'h41F0] = 8'h00;
RAM[16'h41F1] = 8'h00;
RAM[16'h41F2] = 8'h00;
RAM[16'h41F3] = 8'h00;
RAM[16'h41F4] = 8'h00;
RAM[16'h41F5] = 8'h00;
RAM[16'h41F6] = 8'h00;
RAM[16'h41F7] = 8'h00;
RAM[16'h41F8] = 8'h00;
RAM[16'h41F9] = 8'h00;
RAM[16'h41FA] = 8'h00;
RAM[16'h41FB] = 8'h00;
RAM[16'h41FC] = 8'h00;
RAM[16'h41FD] = 8'h00;
RAM[16'h41FE] = 8'h00;
RAM[16'h41FF] = 8'h00;
RAM[16'h4200] = 8'h00;
RAM[16'h4201] = 8'h00;
RAM[16'h4202] = 8'h00;
RAM[16'h4203] = 8'h00;
RAM[16'h4204] = 8'h00;
RAM[16'h4205] = 8'h00;
RAM[16'h4206] = 8'h00;
RAM[16'h4207] = 8'h00;
RAM[16'h4208] = 8'h00;
RAM[16'h4209] = 8'h00;
RAM[16'h420A] = 8'h00;
RAM[16'h420B] = 8'h00;
RAM[16'h420C] = 8'h00;
RAM[16'h420D] = 8'h00;
RAM[16'h420E] = 8'h00;
RAM[16'h420F] = 8'h00;
RAM[16'h4210] = 8'h00;
RAM[16'h4211] = 8'h00;
RAM[16'h4212] = 8'h00;
RAM[16'h4213] = 8'h00;
RAM[16'h4214] = 8'h00;
RAM[16'h4215] = 8'h00;
RAM[16'h4216] = 8'h00;
RAM[16'h4217] = 8'h00;
RAM[16'h4218] = 8'h00;
RAM[16'h4219] = 8'h00;
RAM[16'h421A] = 8'h00;
RAM[16'h421B] = 8'h00;
RAM[16'h421C] = 8'h00;
RAM[16'h421D] = 8'h00;
RAM[16'h421E] = 8'h00;
RAM[16'h421F] = 8'h00;
RAM[16'h4220] = 8'h00;
RAM[16'h4221] = 8'h00;
RAM[16'h4222] = 8'h00;
RAM[16'h4223] = 8'h00;
RAM[16'h4224] = 8'h00;
RAM[16'h4225] = 8'h00;
RAM[16'h4226] = 8'h00;
RAM[16'h4227] = 8'h00;
RAM[16'h4228] = 8'h00;
RAM[16'h4229] = 8'h00;
RAM[16'h422A] = 8'h00;
RAM[16'h422B] = 8'h00;
RAM[16'h422C] = 8'h00;
RAM[16'h422D] = 8'h00;
RAM[16'h422E] = 8'h00;
RAM[16'h422F] = 8'h00;
RAM[16'h4230] = 8'h00;
RAM[16'h4231] = 8'h00;
RAM[16'h4232] = 8'h00;
RAM[16'h4233] = 8'h00;
RAM[16'h4234] = 8'h00;
RAM[16'h4235] = 8'h00;
RAM[16'h4236] = 8'h00;
RAM[16'h4237] = 8'h00;
RAM[16'h4238] = 8'h00;
RAM[16'h4239] = 8'h00;
RAM[16'h423A] = 8'h00;
RAM[16'h423B] = 8'h00;
RAM[16'h423C] = 8'h00;
RAM[16'h423D] = 8'h00;
RAM[16'h423E] = 8'h00;
RAM[16'h423F] = 8'h00;
RAM[16'h4240] = 8'h00;
RAM[16'h4241] = 8'h00;
RAM[16'h4242] = 8'h00;
RAM[16'h4243] = 8'h00;
RAM[16'h4244] = 8'h00;
RAM[16'h4245] = 8'h00;
RAM[16'h4246] = 8'h00;
RAM[16'h4247] = 8'h00;
RAM[16'h4248] = 8'h00;
RAM[16'h4249] = 8'h00;
RAM[16'h424A] = 8'h00;
RAM[16'h424B] = 8'h00;
RAM[16'h424C] = 8'h00;
RAM[16'h424D] = 8'h00;
RAM[16'h424E] = 8'h00;
RAM[16'h424F] = 8'h00;
RAM[16'h4250] = 8'h00;
RAM[16'h4251] = 8'h00;
RAM[16'h4252] = 8'h00;
RAM[16'h4253] = 8'h00;
RAM[16'h4254] = 8'h00;
RAM[16'h4255] = 8'h00;
RAM[16'h4256] = 8'h00;
RAM[16'h4257] = 8'h00;
RAM[16'h4258] = 8'h00;
RAM[16'h4259] = 8'h00;
RAM[16'h425A] = 8'h00;
RAM[16'h425B] = 8'h00;
RAM[16'h425C] = 8'h00;
RAM[16'h425D] = 8'h00;
RAM[16'h425E] = 8'h00;
RAM[16'h425F] = 8'h00;
RAM[16'h4260] = 8'h00;
RAM[16'h4261] = 8'h00;
RAM[16'h4262] = 8'h00;
RAM[16'h4263] = 8'h00;
RAM[16'h4264] = 8'h00;
RAM[16'h4265] = 8'h00;
RAM[16'h4266] = 8'h00;
RAM[16'h4267] = 8'h00;
RAM[16'h4268] = 8'h00;
RAM[16'h4269] = 8'h00;
RAM[16'h426A] = 8'h00;
RAM[16'h426B] = 8'h00;
RAM[16'h426C] = 8'h00;
RAM[16'h426D] = 8'h00;
RAM[16'h426E] = 8'h00;
RAM[16'h426F] = 8'h00;
RAM[16'h4270] = 8'h00;
RAM[16'h4271] = 8'h00;
RAM[16'h4272] = 8'h00;
RAM[16'h4273] = 8'h00;
RAM[16'h4274] = 8'h00;
RAM[16'h4275] = 8'h00;
RAM[16'h4276] = 8'h00;
RAM[16'h4277] = 8'h00;
RAM[16'h4278] = 8'h00;
RAM[16'h4279] = 8'h00;
RAM[16'h427A] = 8'h00;
RAM[16'h427B] = 8'h00;
RAM[16'h427C] = 8'h00;
RAM[16'h427D] = 8'h00;
RAM[16'h427E] = 8'h00;
RAM[16'h427F] = 8'h00;
RAM[16'h4280] = 8'h00;
RAM[16'h4281] = 8'h00;
RAM[16'h4282] = 8'h00;
RAM[16'h4283] = 8'h00;
RAM[16'h4284] = 8'h00;
RAM[16'h4285] = 8'h00;
RAM[16'h4286] = 8'h00;
RAM[16'h4287] = 8'h00;
RAM[16'h4288] = 8'h00;
RAM[16'h4289] = 8'h00;
RAM[16'h428A] = 8'h00;
RAM[16'h428B] = 8'h00;
RAM[16'h428C] = 8'h00;
RAM[16'h428D] = 8'h00;
RAM[16'h428E] = 8'h00;
RAM[16'h428F] = 8'h00;
RAM[16'h4290] = 8'h00;
RAM[16'h4291] = 8'h00;
RAM[16'h4292] = 8'h00;
RAM[16'h4293] = 8'h00;
RAM[16'h4294] = 8'h00;
RAM[16'h4295] = 8'h00;
RAM[16'h4296] = 8'h00;
RAM[16'h4297] = 8'h00;
RAM[16'h4298] = 8'h00;
RAM[16'h4299] = 8'h00;
RAM[16'h429A] = 8'h00;
RAM[16'h429B] = 8'h00;
RAM[16'h429C] = 8'h00;
RAM[16'h429D] = 8'h00;
RAM[16'h429E] = 8'h00;
RAM[16'h429F] = 8'h00;
RAM[16'h42A0] = 8'h00;
RAM[16'h42A1] = 8'h00;
RAM[16'h42A2] = 8'h00;
RAM[16'h42A3] = 8'h00;
RAM[16'h42A4] = 8'h00;
RAM[16'h42A5] = 8'h00;
RAM[16'h42A6] = 8'h00;
RAM[16'h42A7] = 8'h00;
RAM[16'h42A8] = 8'h00;
RAM[16'h42A9] = 8'h00;
RAM[16'h42AA] = 8'h00;
RAM[16'h42AB] = 8'h00;
RAM[16'h42AC] = 8'h00;
RAM[16'h42AD] = 8'h00;
RAM[16'h42AE] = 8'h00;
RAM[16'h42AF] = 8'h00;
RAM[16'h42B0] = 8'h00;
RAM[16'h42B1] = 8'h00;
RAM[16'h42B2] = 8'h00;
RAM[16'h42B3] = 8'h00;
RAM[16'h42B4] = 8'h00;
RAM[16'h42B5] = 8'h00;
RAM[16'h42B6] = 8'h00;
RAM[16'h42B7] = 8'h00;
RAM[16'h42B8] = 8'h00;
RAM[16'h42B9] = 8'h00;
RAM[16'h42BA] = 8'h00;
RAM[16'h42BB] = 8'h00;
RAM[16'h42BC] = 8'h00;
RAM[16'h42BD] = 8'h00;
RAM[16'h42BE] = 8'h00;
RAM[16'h42BF] = 8'h00;
RAM[16'h42C0] = 8'h00;
RAM[16'h42C1] = 8'h00;
RAM[16'h42C2] = 8'h00;
RAM[16'h42C3] = 8'h00;
RAM[16'h42C4] = 8'h00;
RAM[16'h42C5] = 8'h00;
RAM[16'h42C6] = 8'h00;
RAM[16'h42C7] = 8'h00;
RAM[16'h42C8] = 8'h00;
RAM[16'h42C9] = 8'h00;
RAM[16'h42CA] = 8'h00;
RAM[16'h42CB] = 8'h00;
RAM[16'h42CC] = 8'h00;
RAM[16'h42CD] = 8'h00;
RAM[16'h42CE] = 8'h00;
RAM[16'h42CF] = 8'h00;
RAM[16'h42D0] = 8'h00;
RAM[16'h42D1] = 8'h00;
RAM[16'h42D2] = 8'h00;
RAM[16'h42D3] = 8'h00;
RAM[16'h42D4] = 8'h00;
RAM[16'h42D5] = 8'h00;
RAM[16'h42D6] = 8'h00;
RAM[16'h42D7] = 8'h00;
RAM[16'h42D8] = 8'h00;
RAM[16'h42D9] = 8'h00;
RAM[16'h42DA] = 8'h00;
RAM[16'h42DB] = 8'h00;
RAM[16'h42DC] = 8'h00;
RAM[16'h42DD] = 8'h00;
RAM[16'h42DE] = 8'h00;
RAM[16'h42DF] = 8'h00;
RAM[16'h42E0] = 8'h00;
RAM[16'h42E1] = 8'h00;
RAM[16'h42E2] = 8'h00;
RAM[16'h42E3] = 8'h00;
RAM[16'h42E4] = 8'h00;
RAM[16'h42E5] = 8'h00;
RAM[16'h42E6] = 8'h00;
RAM[16'h42E7] = 8'h00;
RAM[16'h42E8] = 8'h00;
RAM[16'h42E9] = 8'h00;
RAM[16'h42EA] = 8'h00;
RAM[16'h42EB] = 8'h00;
RAM[16'h42EC] = 8'h00;
RAM[16'h42ED] = 8'h00;
RAM[16'h42EE] = 8'h00;
RAM[16'h42EF] = 8'h00;
RAM[16'h42F0] = 8'h00;
RAM[16'h42F1] = 8'h00;
RAM[16'h42F2] = 8'h00;
RAM[16'h42F3] = 8'h00;
RAM[16'h42F4] = 8'h00;
RAM[16'h42F5] = 8'h00;
RAM[16'h42F6] = 8'h00;
RAM[16'h42F7] = 8'h00;
RAM[16'h42F8] = 8'h00;
RAM[16'h42F9] = 8'h00;
RAM[16'h42FA] = 8'h00;
RAM[16'h42FB] = 8'h00;
RAM[16'h42FC] = 8'h00;
RAM[16'h42FD] = 8'h00;
RAM[16'h42FE] = 8'h00;
RAM[16'h42FF] = 8'h00;
RAM[16'h4300] = 8'h00;
RAM[16'h4301] = 8'h00;
RAM[16'h4302] = 8'h00;
RAM[16'h4303] = 8'h00;
RAM[16'h4304] = 8'h00;
RAM[16'h4305] = 8'h00;
RAM[16'h4306] = 8'h00;
RAM[16'h4307] = 8'h00;
RAM[16'h4308] = 8'h00;
RAM[16'h4309] = 8'h00;
RAM[16'h430A] = 8'h00;
RAM[16'h430B] = 8'h00;
RAM[16'h430C] = 8'h00;
RAM[16'h430D] = 8'h00;
RAM[16'h430E] = 8'h00;
RAM[16'h430F] = 8'h00;
RAM[16'h4310] = 8'h00;
RAM[16'h4311] = 8'h00;
RAM[16'h4312] = 8'h00;
RAM[16'h4313] = 8'h00;
RAM[16'h4314] = 8'h00;
RAM[16'h4315] = 8'h00;
RAM[16'h4316] = 8'h00;
RAM[16'h4317] = 8'h00;
RAM[16'h4318] = 8'h00;
RAM[16'h4319] = 8'h00;
RAM[16'h431A] = 8'h00;
RAM[16'h431B] = 8'h00;
RAM[16'h431C] = 8'h00;
RAM[16'h431D] = 8'h00;
RAM[16'h431E] = 8'h00;
RAM[16'h431F] = 8'h00;
RAM[16'h4320] = 8'h00;
RAM[16'h4321] = 8'h00;
RAM[16'h4322] = 8'h00;
RAM[16'h4323] = 8'h00;
RAM[16'h4324] = 8'h00;
RAM[16'h4325] = 8'h00;
RAM[16'h4326] = 8'h00;
RAM[16'h4327] = 8'h00;
RAM[16'h4328] = 8'h00;
RAM[16'h4329] = 8'h00;
RAM[16'h432A] = 8'h00;
RAM[16'h432B] = 8'h00;
RAM[16'h432C] = 8'h00;
RAM[16'h432D] = 8'h00;
RAM[16'h432E] = 8'h00;
RAM[16'h432F] = 8'h00;
RAM[16'h4330] = 8'h00;
RAM[16'h4331] = 8'h00;
RAM[16'h4332] = 8'h00;
RAM[16'h4333] = 8'h00;
RAM[16'h4334] = 8'h00;
RAM[16'h4335] = 8'h00;
RAM[16'h4336] = 8'h00;
RAM[16'h4337] = 8'h00;
RAM[16'h4338] = 8'h00;
RAM[16'h4339] = 8'h00;
RAM[16'h433A] = 8'h00;
RAM[16'h433B] = 8'h00;
RAM[16'h433C] = 8'h00;
RAM[16'h433D] = 8'h00;
RAM[16'h433E] = 8'h00;
RAM[16'h433F] = 8'h00;
RAM[16'h4340] = 8'h00;
RAM[16'h4341] = 8'h00;
RAM[16'h4342] = 8'h00;
RAM[16'h4343] = 8'h00;
RAM[16'h4344] = 8'h00;
RAM[16'h4345] = 8'h00;
RAM[16'h4346] = 8'h00;
RAM[16'h4347] = 8'h00;
RAM[16'h4348] = 8'h00;
RAM[16'h4349] = 8'h00;
RAM[16'h434A] = 8'h00;
RAM[16'h434B] = 8'h00;
RAM[16'h434C] = 8'h00;
RAM[16'h434D] = 8'h00;
RAM[16'h434E] = 8'h00;
RAM[16'h434F] = 8'h00;
RAM[16'h4350] = 8'h00;
RAM[16'h4351] = 8'h00;
RAM[16'h4352] = 8'h00;
RAM[16'h4353] = 8'h00;
RAM[16'h4354] = 8'h00;
RAM[16'h4355] = 8'h00;
RAM[16'h4356] = 8'h00;
RAM[16'h4357] = 8'h00;
RAM[16'h4358] = 8'h00;
RAM[16'h4359] = 8'h00;
RAM[16'h435A] = 8'h00;
RAM[16'h435B] = 8'h00;
RAM[16'h435C] = 8'h00;
RAM[16'h435D] = 8'h00;
RAM[16'h435E] = 8'h00;
RAM[16'h435F] = 8'h00;
RAM[16'h4360] = 8'h00;
RAM[16'h4361] = 8'h00;
RAM[16'h4362] = 8'h00;
RAM[16'h4363] = 8'h00;
RAM[16'h4364] = 8'h00;
RAM[16'h4365] = 8'h00;
RAM[16'h4366] = 8'h00;
RAM[16'h4367] = 8'h00;
RAM[16'h4368] = 8'h00;
RAM[16'h4369] = 8'h00;
RAM[16'h436A] = 8'h00;
RAM[16'h436B] = 8'h00;
RAM[16'h436C] = 8'h00;
RAM[16'h436D] = 8'h00;
RAM[16'h436E] = 8'h00;
RAM[16'h436F] = 8'h00;
RAM[16'h4370] = 8'h00;
RAM[16'h4371] = 8'h00;
RAM[16'h4372] = 8'h00;
RAM[16'h4373] = 8'h00;
RAM[16'h4374] = 8'h00;
RAM[16'h4375] = 8'h00;
RAM[16'h4376] = 8'h00;
RAM[16'h4377] = 8'h00;
RAM[16'h4378] = 8'h00;
RAM[16'h4379] = 8'h00;
RAM[16'h437A] = 8'h00;
RAM[16'h437B] = 8'h00;
RAM[16'h437C] = 8'h00;
RAM[16'h437D] = 8'h00;
RAM[16'h437E] = 8'h00;
RAM[16'h437F] = 8'h00;
RAM[16'h4380] = 8'h00;
RAM[16'h4381] = 8'h00;
RAM[16'h4382] = 8'h00;
RAM[16'h4383] = 8'h00;
RAM[16'h4384] = 8'h00;
RAM[16'h4385] = 8'h00;
RAM[16'h4386] = 8'h00;
RAM[16'h4387] = 8'h00;
RAM[16'h4388] = 8'h00;
RAM[16'h4389] = 8'h00;
RAM[16'h438A] = 8'h00;
RAM[16'h438B] = 8'h00;
RAM[16'h438C] = 8'h00;
RAM[16'h438D] = 8'h00;
RAM[16'h438E] = 8'h00;
RAM[16'h438F] = 8'h00;
RAM[16'h4390] = 8'h00;
RAM[16'h4391] = 8'h00;
RAM[16'h4392] = 8'h00;
RAM[16'h4393] = 8'h00;
RAM[16'h4394] = 8'h00;
RAM[16'h4395] = 8'h00;
RAM[16'h4396] = 8'h00;
RAM[16'h4397] = 8'h00;
RAM[16'h4398] = 8'h00;
RAM[16'h4399] = 8'h00;
RAM[16'h439A] = 8'h00;
RAM[16'h439B] = 8'h00;
RAM[16'h439C] = 8'h00;
RAM[16'h439D] = 8'h00;
RAM[16'h439E] = 8'h00;
RAM[16'h439F] = 8'h00;
RAM[16'h43A0] = 8'h00;
RAM[16'h43A1] = 8'h00;
RAM[16'h43A2] = 8'h00;
RAM[16'h43A3] = 8'h00;
RAM[16'h43A4] = 8'h00;
RAM[16'h43A5] = 8'h00;
RAM[16'h43A6] = 8'h00;
RAM[16'h43A7] = 8'h00;
RAM[16'h43A8] = 8'h00;
RAM[16'h43A9] = 8'h00;
RAM[16'h43AA] = 8'h00;
RAM[16'h43AB] = 8'h00;
RAM[16'h43AC] = 8'h00;
RAM[16'h43AD] = 8'h00;
RAM[16'h43AE] = 8'h00;
RAM[16'h43AF] = 8'h00;
RAM[16'h43B0] = 8'h00;
RAM[16'h43B1] = 8'h00;
RAM[16'h43B2] = 8'h00;
RAM[16'h43B3] = 8'h00;
RAM[16'h43B4] = 8'h00;
RAM[16'h43B5] = 8'h00;
RAM[16'h43B6] = 8'h00;
RAM[16'h43B7] = 8'h00;
RAM[16'h43B8] = 8'h00;
RAM[16'h43B9] = 8'h00;
RAM[16'h43BA] = 8'h00;
RAM[16'h43BB] = 8'h00;
RAM[16'h43BC] = 8'h00;
RAM[16'h43BD] = 8'h00;
RAM[16'h43BE] = 8'h00;
RAM[16'h43BF] = 8'h00;
RAM[16'h43C0] = 8'h00;
RAM[16'h43C1] = 8'h00;
RAM[16'h43C2] = 8'h00;
RAM[16'h43C3] = 8'h00;
RAM[16'h43C4] = 8'h00;
RAM[16'h43C5] = 8'h00;
RAM[16'h43C6] = 8'h00;
RAM[16'h43C7] = 8'h00;
RAM[16'h43C8] = 8'h00;
RAM[16'h43C9] = 8'h00;
RAM[16'h43CA] = 8'h00;
RAM[16'h43CB] = 8'h00;
RAM[16'h43CC] = 8'h00;
RAM[16'h43CD] = 8'h00;
RAM[16'h43CE] = 8'h00;
RAM[16'h43CF] = 8'h00;
RAM[16'h43D0] = 8'h00;
RAM[16'h43D1] = 8'h00;
RAM[16'h43D2] = 8'h00;
RAM[16'h43D3] = 8'h00;
RAM[16'h43D4] = 8'h00;
RAM[16'h43D5] = 8'h00;
RAM[16'h43D6] = 8'h00;
RAM[16'h43D7] = 8'h00;
RAM[16'h43D8] = 8'h00;
RAM[16'h43D9] = 8'h00;
RAM[16'h43DA] = 8'h00;
RAM[16'h43DB] = 8'h00;
RAM[16'h43DC] = 8'h00;
RAM[16'h43DD] = 8'h00;
RAM[16'h43DE] = 8'h00;
RAM[16'h43DF] = 8'h00;
RAM[16'h43E0] = 8'h00;
RAM[16'h43E1] = 8'h00;
RAM[16'h43E2] = 8'h00;
RAM[16'h43E3] = 8'h00;
RAM[16'h43E4] = 8'h00;
RAM[16'h43E5] = 8'h00;
RAM[16'h43E6] = 8'h00;
RAM[16'h43E7] = 8'h00;
RAM[16'h43E8] = 8'h00;
RAM[16'h43E9] = 8'h00;
RAM[16'h43EA] = 8'h00;
RAM[16'h43EB] = 8'h00;
RAM[16'h43EC] = 8'h00;
RAM[16'h43ED] = 8'h00;
RAM[16'h43EE] = 8'h00;
RAM[16'h43EF] = 8'h00;
RAM[16'h43F0] = 8'h00;
RAM[16'h43F1] = 8'h00;
RAM[16'h43F2] = 8'h00;
RAM[16'h43F3] = 8'h00;
RAM[16'h43F4] = 8'h00;
RAM[16'h43F5] = 8'h00;
RAM[16'h43F6] = 8'h00;
RAM[16'h43F7] = 8'h00;
RAM[16'h43F8] = 8'h00;
RAM[16'h43F9] = 8'h00;
RAM[16'h43FA] = 8'h00;
RAM[16'h43FB] = 8'h00;
RAM[16'h43FC] = 8'h00;
RAM[16'h43FD] = 8'h00;
RAM[16'h43FE] = 8'h00;
RAM[16'h43FF] = 8'h00;
RAM[16'h4400] = 8'h00;
RAM[16'h4401] = 8'h00;
RAM[16'h4402] = 8'h00;
RAM[16'h4403] = 8'h00;
RAM[16'h4404] = 8'h00;
RAM[16'h4405] = 8'h00;
RAM[16'h4406] = 8'h00;
RAM[16'h4407] = 8'h00;
RAM[16'h4408] = 8'h00;
RAM[16'h4409] = 8'h00;
RAM[16'h440A] = 8'h00;
RAM[16'h440B] = 8'h00;
RAM[16'h440C] = 8'h00;
RAM[16'h440D] = 8'h00;
RAM[16'h440E] = 8'h00;
RAM[16'h440F] = 8'h00;
RAM[16'h4410] = 8'h00;
RAM[16'h4411] = 8'h00;
RAM[16'h4412] = 8'h00;
RAM[16'h4413] = 8'h00;
RAM[16'h4414] = 8'h00;
RAM[16'h4415] = 8'h00;
RAM[16'h4416] = 8'h00;
RAM[16'h4417] = 8'h00;
RAM[16'h4418] = 8'h00;
RAM[16'h4419] = 8'h00;
RAM[16'h441A] = 8'h00;
RAM[16'h441B] = 8'h00;
RAM[16'h441C] = 8'h00;
RAM[16'h441D] = 8'h00;
RAM[16'h441E] = 8'h00;
RAM[16'h441F] = 8'h00;
RAM[16'h4420] = 8'h00;
RAM[16'h4421] = 8'h00;
RAM[16'h4422] = 8'h00;
RAM[16'h4423] = 8'h00;
RAM[16'h4424] = 8'h00;
RAM[16'h4425] = 8'h00;
RAM[16'h4426] = 8'h00;
RAM[16'h4427] = 8'h00;
RAM[16'h4428] = 8'h00;
RAM[16'h4429] = 8'h00;
RAM[16'h442A] = 8'h00;
RAM[16'h442B] = 8'h00;
RAM[16'h442C] = 8'h00;
RAM[16'h442D] = 8'h00;
RAM[16'h442E] = 8'h00;
RAM[16'h442F] = 8'h00;
RAM[16'h4430] = 8'h00;
RAM[16'h4431] = 8'h00;
RAM[16'h4432] = 8'h00;
RAM[16'h4433] = 8'h00;
RAM[16'h4434] = 8'h00;
RAM[16'h4435] = 8'h00;
RAM[16'h4436] = 8'h00;
RAM[16'h4437] = 8'h00;
RAM[16'h4438] = 8'h00;
RAM[16'h4439] = 8'h00;
RAM[16'h443A] = 8'h00;
RAM[16'h443B] = 8'h00;
RAM[16'h443C] = 8'h00;
RAM[16'h443D] = 8'h00;
RAM[16'h443E] = 8'h00;
RAM[16'h443F] = 8'h00;
RAM[16'h4440] = 8'h00;
RAM[16'h4441] = 8'h00;
RAM[16'h4442] = 8'h00;
RAM[16'h4443] = 8'h00;
RAM[16'h4444] = 8'h00;
RAM[16'h4445] = 8'h00;
RAM[16'h4446] = 8'h00;
RAM[16'h4447] = 8'h00;
RAM[16'h4448] = 8'h00;
RAM[16'h4449] = 8'h00;
RAM[16'h444A] = 8'h00;
RAM[16'h444B] = 8'h00;
RAM[16'h444C] = 8'h00;
RAM[16'h444D] = 8'h00;
RAM[16'h444E] = 8'h00;
RAM[16'h444F] = 8'h00;
RAM[16'h4450] = 8'h00;
RAM[16'h4451] = 8'h00;
RAM[16'h4452] = 8'h00;
RAM[16'h4453] = 8'h00;
RAM[16'h4454] = 8'h00;
RAM[16'h4455] = 8'h00;
RAM[16'h4456] = 8'h00;
RAM[16'h4457] = 8'h00;
RAM[16'h4458] = 8'h00;
RAM[16'h4459] = 8'h00;
RAM[16'h445A] = 8'h00;
RAM[16'h445B] = 8'h00;
RAM[16'h445C] = 8'h00;
RAM[16'h445D] = 8'h00;
RAM[16'h445E] = 8'h00;
RAM[16'h445F] = 8'h00;
RAM[16'h4460] = 8'h00;
RAM[16'h4461] = 8'h00;
RAM[16'h4462] = 8'h00;
RAM[16'h4463] = 8'h00;
RAM[16'h4464] = 8'h00;
RAM[16'h4465] = 8'h00;
RAM[16'h4466] = 8'h00;
RAM[16'h4467] = 8'h00;
RAM[16'h4468] = 8'h00;
RAM[16'h4469] = 8'h00;
RAM[16'h446A] = 8'h00;
RAM[16'h446B] = 8'h00;
RAM[16'h446C] = 8'h00;
RAM[16'h446D] = 8'h00;
RAM[16'h446E] = 8'h00;
RAM[16'h446F] = 8'h00;
RAM[16'h4470] = 8'h00;
RAM[16'h4471] = 8'h00;
RAM[16'h4472] = 8'h00;
RAM[16'h4473] = 8'h00;
RAM[16'h4474] = 8'h00;
RAM[16'h4475] = 8'h00;
RAM[16'h4476] = 8'h00;
RAM[16'h4477] = 8'h00;
RAM[16'h4478] = 8'h00;
RAM[16'h4479] = 8'h00;
RAM[16'h447A] = 8'h00;
RAM[16'h447B] = 8'h00;
RAM[16'h447C] = 8'h00;
RAM[16'h447D] = 8'h00;
RAM[16'h447E] = 8'h00;
RAM[16'h447F] = 8'h00;
RAM[16'h4480] = 8'h00;
RAM[16'h4481] = 8'h00;
RAM[16'h4482] = 8'h00;
RAM[16'h4483] = 8'h00;
RAM[16'h4484] = 8'h00;
RAM[16'h4485] = 8'h00;
RAM[16'h4486] = 8'h00;
RAM[16'h4487] = 8'h00;
RAM[16'h4488] = 8'h00;
RAM[16'h4489] = 8'h00;
RAM[16'h448A] = 8'h00;
RAM[16'h448B] = 8'h00;
RAM[16'h448C] = 8'h00;
RAM[16'h448D] = 8'h00;
RAM[16'h448E] = 8'h00;
RAM[16'h448F] = 8'h00;
RAM[16'h4490] = 8'h00;
RAM[16'h4491] = 8'h00;
RAM[16'h4492] = 8'h00;
RAM[16'h4493] = 8'h00;
RAM[16'h4494] = 8'h00;
RAM[16'h4495] = 8'h00;
RAM[16'h4496] = 8'h00;
RAM[16'h4497] = 8'h00;
RAM[16'h4498] = 8'h00;
RAM[16'h4499] = 8'h00;
RAM[16'h449A] = 8'h00;
RAM[16'h449B] = 8'h00;
RAM[16'h449C] = 8'h00;
RAM[16'h449D] = 8'h00;
RAM[16'h449E] = 8'h00;
RAM[16'h449F] = 8'h00;
RAM[16'h44A0] = 8'h00;
RAM[16'h44A1] = 8'h00;
RAM[16'h44A2] = 8'h00;
RAM[16'h44A3] = 8'h00;
RAM[16'h44A4] = 8'h00;
RAM[16'h44A5] = 8'h00;
RAM[16'h44A6] = 8'h00;
RAM[16'h44A7] = 8'h00;
RAM[16'h44A8] = 8'h00;
RAM[16'h44A9] = 8'h00;
RAM[16'h44AA] = 8'h00;
RAM[16'h44AB] = 8'h00;
RAM[16'h44AC] = 8'h00;
RAM[16'h44AD] = 8'h00;
RAM[16'h44AE] = 8'h00;
RAM[16'h44AF] = 8'h00;
RAM[16'h44B0] = 8'h00;
RAM[16'h44B1] = 8'h00;
RAM[16'h44B2] = 8'h00;
RAM[16'h44B3] = 8'h00;
RAM[16'h44B4] = 8'h00;
RAM[16'h44B5] = 8'h00;
RAM[16'h44B6] = 8'h00;
RAM[16'h44B7] = 8'h00;
RAM[16'h44B8] = 8'h00;
RAM[16'h44B9] = 8'h00;
RAM[16'h44BA] = 8'h00;
RAM[16'h44BB] = 8'h00;
RAM[16'h44BC] = 8'h00;
RAM[16'h44BD] = 8'h00;
RAM[16'h44BE] = 8'h00;
RAM[16'h44BF] = 8'h00;
RAM[16'h44C0] = 8'h00;
RAM[16'h44C1] = 8'h00;
RAM[16'h44C2] = 8'h00;
RAM[16'h44C3] = 8'h00;
RAM[16'h44C4] = 8'h00;
RAM[16'h44C5] = 8'h00;
RAM[16'h44C6] = 8'h00;
RAM[16'h44C7] = 8'h00;
RAM[16'h44C8] = 8'h00;
RAM[16'h44C9] = 8'h00;
RAM[16'h44CA] = 8'h00;
RAM[16'h44CB] = 8'h00;
RAM[16'h44CC] = 8'h00;
RAM[16'h44CD] = 8'h00;
RAM[16'h44CE] = 8'h00;
RAM[16'h44CF] = 8'h00;
RAM[16'h44D0] = 8'h00;
RAM[16'h44D1] = 8'h00;
RAM[16'h44D2] = 8'h00;
RAM[16'h44D3] = 8'h00;
RAM[16'h44D4] = 8'h00;
RAM[16'h44D5] = 8'h00;
RAM[16'h44D6] = 8'h00;
RAM[16'h44D7] = 8'h00;
RAM[16'h44D8] = 8'h00;
RAM[16'h44D9] = 8'h00;
RAM[16'h44DA] = 8'h00;
RAM[16'h44DB] = 8'h00;
RAM[16'h44DC] = 8'h00;
RAM[16'h44DD] = 8'h00;
RAM[16'h44DE] = 8'h00;
RAM[16'h44DF] = 8'h00;
RAM[16'h44E0] = 8'h00;
RAM[16'h44E1] = 8'h00;
RAM[16'h44E2] = 8'h00;
RAM[16'h44E3] = 8'h00;
RAM[16'h44E4] = 8'h00;
RAM[16'h44E5] = 8'h00;
RAM[16'h44E6] = 8'h00;
RAM[16'h44E7] = 8'h00;
RAM[16'h44E8] = 8'h00;
RAM[16'h44E9] = 8'h00;
RAM[16'h44EA] = 8'h00;
RAM[16'h44EB] = 8'h00;
RAM[16'h44EC] = 8'h00;
RAM[16'h44ED] = 8'h00;
RAM[16'h44EE] = 8'h00;
RAM[16'h44EF] = 8'h00;
RAM[16'h44F0] = 8'h00;
RAM[16'h44F1] = 8'h00;
RAM[16'h44F2] = 8'h00;
RAM[16'h44F3] = 8'h00;
RAM[16'h44F4] = 8'h00;
RAM[16'h44F5] = 8'h00;
RAM[16'h44F6] = 8'h00;
RAM[16'h44F7] = 8'h00;
RAM[16'h44F8] = 8'h00;
RAM[16'h44F9] = 8'h00;
RAM[16'h44FA] = 8'h00;
RAM[16'h44FB] = 8'h00;
RAM[16'h44FC] = 8'h00;
RAM[16'h44FD] = 8'h00;
RAM[16'h44FE] = 8'h00;
RAM[16'h44FF] = 8'h00;
RAM[16'h4500] = 8'h00;
RAM[16'h4501] = 8'h00;
RAM[16'h4502] = 8'h00;
RAM[16'h4503] = 8'h00;
RAM[16'h4504] = 8'h00;
RAM[16'h4505] = 8'h00;
RAM[16'h4506] = 8'h00;
RAM[16'h4507] = 8'h00;
RAM[16'h4508] = 8'h00;
RAM[16'h4509] = 8'h00;
RAM[16'h450A] = 8'h00;
RAM[16'h450B] = 8'h00;
RAM[16'h450C] = 8'h00;
RAM[16'h450D] = 8'h00;
RAM[16'h450E] = 8'h00;
RAM[16'h450F] = 8'h00;
RAM[16'h4510] = 8'h00;
RAM[16'h4511] = 8'h00;
RAM[16'h4512] = 8'h00;
RAM[16'h4513] = 8'h00;
RAM[16'h4514] = 8'h00;
RAM[16'h4515] = 8'h00;
RAM[16'h4516] = 8'h00;
RAM[16'h4517] = 8'h00;
RAM[16'h4518] = 8'h00;
RAM[16'h4519] = 8'h00;
RAM[16'h451A] = 8'h00;
RAM[16'h451B] = 8'h00;
RAM[16'h451C] = 8'h00;
RAM[16'h451D] = 8'h00;
RAM[16'h451E] = 8'h00;
RAM[16'h451F] = 8'h00;
RAM[16'h4520] = 8'h00;
RAM[16'h4521] = 8'h00;
RAM[16'h4522] = 8'h00;
RAM[16'h4523] = 8'h00;
RAM[16'h4524] = 8'h00;
RAM[16'h4525] = 8'h00;
RAM[16'h4526] = 8'h00;
RAM[16'h4527] = 8'h00;
RAM[16'h4528] = 8'h00;
RAM[16'h4529] = 8'h00;
RAM[16'h452A] = 8'h00;
RAM[16'h452B] = 8'h00;
RAM[16'h452C] = 8'h00;
RAM[16'h452D] = 8'h00;
RAM[16'h452E] = 8'h00;
RAM[16'h452F] = 8'h00;
RAM[16'h4530] = 8'h00;
RAM[16'h4531] = 8'h00;
RAM[16'h4532] = 8'h00;
RAM[16'h4533] = 8'h00;
RAM[16'h4534] = 8'h00;
RAM[16'h4535] = 8'h00;
RAM[16'h4536] = 8'h00;
RAM[16'h4537] = 8'h00;
RAM[16'h4538] = 8'h00;
RAM[16'h4539] = 8'h00;
RAM[16'h453A] = 8'h00;
RAM[16'h453B] = 8'h00;
RAM[16'h453C] = 8'h00;
RAM[16'h453D] = 8'h00;
RAM[16'h453E] = 8'h00;
RAM[16'h453F] = 8'h00;
RAM[16'h4540] = 8'h00;
RAM[16'h4541] = 8'h00;
RAM[16'h4542] = 8'h00;
RAM[16'h4543] = 8'h00;
RAM[16'h4544] = 8'h00;
RAM[16'h4545] = 8'h00;
RAM[16'h4546] = 8'h00;
RAM[16'h4547] = 8'h00;
RAM[16'h4548] = 8'h00;
RAM[16'h4549] = 8'h00;
RAM[16'h454A] = 8'h00;
RAM[16'h454B] = 8'h00;
RAM[16'h454C] = 8'h00;
RAM[16'h454D] = 8'h00;
RAM[16'h454E] = 8'h00;
RAM[16'h454F] = 8'h00;
RAM[16'h4550] = 8'h00;
RAM[16'h4551] = 8'h00;
RAM[16'h4552] = 8'h00;
RAM[16'h4553] = 8'h00;
RAM[16'h4554] = 8'h00;
RAM[16'h4555] = 8'h00;
RAM[16'h4556] = 8'h00;
RAM[16'h4557] = 8'h00;
RAM[16'h4558] = 8'h00;
RAM[16'h4559] = 8'h00;
RAM[16'h455A] = 8'h00;
RAM[16'h455B] = 8'h00;
RAM[16'h455C] = 8'h00;
RAM[16'h455D] = 8'h00;
RAM[16'h455E] = 8'h00;
RAM[16'h455F] = 8'h00;
RAM[16'h4560] = 8'h00;
RAM[16'h4561] = 8'h00;
RAM[16'h4562] = 8'h00;
RAM[16'h4563] = 8'h00;
RAM[16'h4564] = 8'h00;
RAM[16'h4565] = 8'h00;
RAM[16'h4566] = 8'h00;
RAM[16'h4567] = 8'h00;
RAM[16'h4568] = 8'h00;
RAM[16'h4569] = 8'h00;
RAM[16'h456A] = 8'h00;
RAM[16'h456B] = 8'h00;
RAM[16'h456C] = 8'h00;
RAM[16'h456D] = 8'h00;
RAM[16'h456E] = 8'h00;
RAM[16'h456F] = 8'h00;
RAM[16'h4570] = 8'h00;
RAM[16'h4571] = 8'h00;
RAM[16'h4572] = 8'h00;
RAM[16'h4573] = 8'h00;
RAM[16'h4574] = 8'h00;
RAM[16'h4575] = 8'h00;
RAM[16'h4576] = 8'h00;
RAM[16'h4577] = 8'h00;
RAM[16'h4578] = 8'h00;
RAM[16'h4579] = 8'h00;
RAM[16'h457A] = 8'h00;
RAM[16'h457B] = 8'h00;
RAM[16'h457C] = 8'h00;
RAM[16'h457D] = 8'h00;
RAM[16'h457E] = 8'h00;
RAM[16'h457F] = 8'h00;
RAM[16'h4580] = 8'h00;
RAM[16'h4581] = 8'h00;
RAM[16'h4582] = 8'h00;
RAM[16'h4583] = 8'h00;
RAM[16'h4584] = 8'h00;
RAM[16'h4585] = 8'h00;
RAM[16'h4586] = 8'h00;
RAM[16'h4587] = 8'h00;
RAM[16'h4588] = 8'h00;
RAM[16'h4589] = 8'h00;
RAM[16'h458A] = 8'h00;
RAM[16'h458B] = 8'h00;
RAM[16'h458C] = 8'h00;
RAM[16'h458D] = 8'h00;
RAM[16'h458E] = 8'h00;
RAM[16'h458F] = 8'h00;
RAM[16'h4590] = 8'h00;
RAM[16'h4591] = 8'h00;
RAM[16'h4592] = 8'h00;
RAM[16'h4593] = 8'h00;
RAM[16'h4594] = 8'h00;
RAM[16'h4595] = 8'h00;
RAM[16'h4596] = 8'h00;
RAM[16'h4597] = 8'h00;
RAM[16'h4598] = 8'h00;
RAM[16'h4599] = 8'h00;
RAM[16'h459A] = 8'h00;
RAM[16'h459B] = 8'h00;
RAM[16'h459C] = 8'h00;
RAM[16'h459D] = 8'h00;
RAM[16'h459E] = 8'h00;
RAM[16'h459F] = 8'h00;
RAM[16'h45A0] = 8'h00;
RAM[16'h45A1] = 8'h00;
RAM[16'h45A2] = 8'h00;
RAM[16'h45A3] = 8'h00;
RAM[16'h45A4] = 8'h00;
RAM[16'h45A5] = 8'h00;
RAM[16'h45A6] = 8'h00;
RAM[16'h45A7] = 8'h00;
RAM[16'h45A8] = 8'h00;
RAM[16'h45A9] = 8'h00;
RAM[16'h45AA] = 8'h00;
RAM[16'h45AB] = 8'h00;
RAM[16'h45AC] = 8'h00;
RAM[16'h45AD] = 8'h00;
RAM[16'h45AE] = 8'h00;
RAM[16'h45AF] = 8'h00;
RAM[16'h45B0] = 8'h00;
RAM[16'h45B1] = 8'h00;
RAM[16'h45B2] = 8'h00;
RAM[16'h45B3] = 8'h00;
RAM[16'h45B4] = 8'h00;
RAM[16'h45B5] = 8'h00;
RAM[16'h45B6] = 8'h00;
RAM[16'h45B7] = 8'h00;
RAM[16'h45B8] = 8'h00;
RAM[16'h45B9] = 8'h00;
RAM[16'h45BA] = 8'h00;
RAM[16'h45BB] = 8'h00;
RAM[16'h45BC] = 8'h00;
RAM[16'h45BD] = 8'h00;
RAM[16'h45BE] = 8'h00;
RAM[16'h45BF] = 8'h00;
RAM[16'h45C0] = 8'h00;
RAM[16'h45C1] = 8'h00;
RAM[16'h45C2] = 8'h00;
RAM[16'h45C3] = 8'h00;
RAM[16'h45C4] = 8'h00;
RAM[16'h45C5] = 8'h00;
RAM[16'h45C6] = 8'h00;
RAM[16'h45C7] = 8'h00;
RAM[16'h45C8] = 8'h00;
RAM[16'h45C9] = 8'h00;
RAM[16'h45CA] = 8'h00;
RAM[16'h45CB] = 8'h00;
RAM[16'h45CC] = 8'h00;
RAM[16'h45CD] = 8'h00;
RAM[16'h45CE] = 8'h00;
RAM[16'h45CF] = 8'h00;
RAM[16'h45D0] = 8'h00;
RAM[16'h45D1] = 8'h00;
RAM[16'h45D2] = 8'h00;
RAM[16'h45D3] = 8'h00;
RAM[16'h45D4] = 8'h00;
RAM[16'h45D5] = 8'h00;
RAM[16'h45D6] = 8'h00;
RAM[16'h45D7] = 8'h00;
RAM[16'h45D8] = 8'h00;
RAM[16'h45D9] = 8'h00;
RAM[16'h45DA] = 8'h00;
RAM[16'h45DB] = 8'h00;
RAM[16'h45DC] = 8'h00;
RAM[16'h45DD] = 8'h00;
RAM[16'h45DE] = 8'h00;
RAM[16'h45DF] = 8'h00;
RAM[16'h45E0] = 8'h00;
RAM[16'h45E1] = 8'h00;
RAM[16'h45E2] = 8'h00;
RAM[16'h45E3] = 8'h00;
RAM[16'h45E4] = 8'h00;
RAM[16'h45E5] = 8'h00;
RAM[16'h45E6] = 8'h00;
RAM[16'h45E7] = 8'h00;
RAM[16'h45E8] = 8'h00;
RAM[16'h45E9] = 8'h00;
RAM[16'h45EA] = 8'h00;
RAM[16'h45EB] = 8'h00;
RAM[16'h45EC] = 8'h00;
RAM[16'h45ED] = 8'h00;
RAM[16'h45EE] = 8'h00;
RAM[16'h45EF] = 8'h00;
RAM[16'h45F0] = 8'h00;
RAM[16'h45F1] = 8'h00;
RAM[16'h45F2] = 8'h00;
RAM[16'h45F3] = 8'h00;
RAM[16'h45F4] = 8'h00;
RAM[16'h45F5] = 8'h00;
RAM[16'h45F6] = 8'h00;
RAM[16'h45F7] = 8'h00;
RAM[16'h45F8] = 8'h00;
RAM[16'h45F9] = 8'h00;
RAM[16'h45FA] = 8'h00;
RAM[16'h45FB] = 8'h00;
RAM[16'h45FC] = 8'h00;
RAM[16'h45FD] = 8'h00;
RAM[16'h45FE] = 8'h00;
RAM[16'h45FF] = 8'h00;
RAM[16'h4600] = 8'h00;
RAM[16'h4601] = 8'h00;
RAM[16'h4602] = 8'h00;
RAM[16'h4603] = 8'h00;
RAM[16'h4604] = 8'h00;
RAM[16'h4605] = 8'h00;
RAM[16'h4606] = 8'h00;
RAM[16'h4607] = 8'h00;
RAM[16'h4608] = 8'h00;
RAM[16'h4609] = 8'h00;
RAM[16'h460A] = 8'h00;
RAM[16'h460B] = 8'h00;
RAM[16'h460C] = 8'h00;
RAM[16'h460D] = 8'h00;
RAM[16'h460E] = 8'h00;
RAM[16'h460F] = 8'h00;
RAM[16'h4610] = 8'h00;
RAM[16'h4611] = 8'h00;
RAM[16'h4612] = 8'h00;
RAM[16'h4613] = 8'h00;
RAM[16'h4614] = 8'h00;
RAM[16'h4615] = 8'h00;
RAM[16'h4616] = 8'h00;
RAM[16'h4617] = 8'h00;
RAM[16'h4618] = 8'h00;
RAM[16'h4619] = 8'h00;
RAM[16'h461A] = 8'h00;
RAM[16'h461B] = 8'h00;
RAM[16'h461C] = 8'h00;
RAM[16'h461D] = 8'h00;
RAM[16'h461E] = 8'h00;
RAM[16'h461F] = 8'h00;
RAM[16'h4620] = 8'h00;
RAM[16'h4621] = 8'h00;
RAM[16'h4622] = 8'h00;
RAM[16'h4623] = 8'h00;
RAM[16'h4624] = 8'h00;
RAM[16'h4625] = 8'h00;
RAM[16'h4626] = 8'h00;
RAM[16'h4627] = 8'h00;
RAM[16'h4628] = 8'h00;
RAM[16'h4629] = 8'h00;
RAM[16'h462A] = 8'h00;
RAM[16'h462B] = 8'h00;
RAM[16'h462C] = 8'h00;
RAM[16'h462D] = 8'h00;
RAM[16'h462E] = 8'h00;
RAM[16'h462F] = 8'h00;
RAM[16'h4630] = 8'h00;
RAM[16'h4631] = 8'h00;
RAM[16'h4632] = 8'h00;
RAM[16'h4633] = 8'h00;
RAM[16'h4634] = 8'h00;
RAM[16'h4635] = 8'h00;
RAM[16'h4636] = 8'h00;
RAM[16'h4637] = 8'h00;
RAM[16'h4638] = 8'h00;
RAM[16'h4639] = 8'h00;
RAM[16'h463A] = 8'h00;
RAM[16'h463B] = 8'h00;
RAM[16'h463C] = 8'h00;
RAM[16'h463D] = 8'h00;
RAM[16'h463E] = 8'h00;
RAM[16'h463F] = 8'h00;
RAM[16'h4640] = 8'h00;
RAM[16'h4641] = 8'h00;
RAM[16'h4642] = 8'h00;
RAM[16'h4643] = 8'h00;
RAM[16'h4644] = 8'h00;
RAM[16'h4645] = 8'h00;
RAM[16'h4646] = 8'h00;
RAM[16'h4647] = 8'h00;
RAM[16'h4648] = 8'h00;
RAM[16'h4649] = 8'h00;
RAM[16'h464A] = 8'h00;
RAM[16'h464B] = 8'h00;
RAM[16'h464C] = 8'h00;
RAM[16'h464D] = 8'h00;
RAM[16'h464E] = 8'h00;
RAM[16'h464F] = 8'h00;
RAM[16'h4650] = 8'h00;
RAM[16'h4651] = 8'h00;
RAM[16'h4652] = 8'h00;
RAM[16'h4653] = 8'h00;
RAM[16'h4654] = 8'h00;
RAM[16'h4655] = 8'h00;
RAM[16'h4656] = 8'h00;
RAM[16'h4657] = 8'h00;
RAM[16'h4658] = 8'h00;
RAM[16'h4659] = 8'h00;
RAM[16'h465A] = 8'h00;
RAM[16'h465B] = 8'h00;
RAM[16'h465C] = 8'h00;
RAM[16'h465D] = 8'h00;
RAM[16'h465E] = 8'h00;
RAM[16'h465F] = 8'h00;
RAM[16'h4660] = 8'h00;
RAM[16'h4661] = 8'h00;
RAM[16'h4662] = 8'h00;
RAM[16'h4663] = 8'h00;
RAM[16'h4664] = 8'h00;
RAM[16'h4665] = 8'h00;
RAM[16'h4666] = 8'h00;
RAM[16'h4667] = 8'h00;
RAM[16'h4668] = 8'h00;
RAM[16'h4669] = 8'h00;
RAM[16'h466A] = 8'h00;
RAM[16'h466B] = 8'h00;
RAM[16'h466C] = 8'h00;
RAM[16'h466D] = 8'h00;
RAM[16'h466E] = 8'h00;
RAM[16'h466F] = 8'h00;
RAM[16'h4670] = 8'h00;
RAM[16'h4671] = 8'h00;
RAM[16'h4672] = 8'h00;
RAM[16'h4673] = 8'h00;
RAM[16'h4674] = 8'h00;
RAM[16'h4675] = 8'h00;
RAM[16'h4676] = 8'h00;
RAM[16'h4677] = 8'h00;
RAM[16'h4678] = 8'h00;
RAM[16'h4679] = 8'h00;
RAM[16'h467A] = 8'h00;
RAM[16'h467B] = 8'h00;
RAM[16'h467C] = 8'h00;
RAM[16'h467D] = 8'h00;
RAM[16'h467E] = 8'h00;
RAM[16'h467F] = 8'h00;
RAM[16'h4680] = 8'h00;
RAM[16'h4681] = 8'h00;
RAM[16'h4682] = 8'h00;
RAM[16'h4683] = 8'h00;
RAM[16'h4684] = 8'h00;
RAM[16'h4685] = 8'h00;
RAM[16'h4686] = 8'h00;
RAM[16'h4687] = 8'h00;
RAM[16'h4688] = 8'h00;
RAM[16'h4689] = 8'h00;
RAM[16'h468A] = 8'h00;
RAM[16'h468B] = 8'h00;
RAM[16'h468C] = 8'h00;
RAM[16'h468D] = 8'h00;
RAM[16'h468E] = 8'h00;
RAM[16'h468F] = 8'h00;
RAM[16'h4690] = 8'h00;
RAM[16'h4691] = 8'h00;
RAM[16'h4692] = 8'h00;
RAM[16'h4693] = 8'h00;
RAM[16'h4694] = 8'h00;
RAM[16'h4695] = 8'h00;
RAM[16'h4696] = 8'h00;
RAM[16'h4697] = 8'h00;
RAM[16'h4698] = 8'h00;
RAM[16'h4699] = 8'h00;
RAM[16'h469A] = 8'h00;
RAM[16'h469B] = 8'h00;
RAM[16'h469C] = 8'h00;
RAM[16'h469D] = 8'h00;
RAM[16'h469E] = 8'h00;
RAM[16'h469F] = 8'h00;
RAM[16'h46A0] = 8'h00;
RAM[16'h46A1] = 8'h00;
RAM[16'h46A2] = 8'h00;
RAM[16'h46A3] = 8'h00;
RAM[16'h46A4] = 8'h00;
RAM[16'h46A5] = 8'h00;
RAM[16'h46A6] = 8'h00;
RAM[16'h46A7] = 8'h00;
RAM[16'h46A8] = 8'h00;
RAM[16'h46A9] = 8'h00;
RAM[16'h46AA] = 8'h00;
RAM[16'h46AB] = 8'h00;
RAM[16'h46AC] = 8'h00;
RAM[16'h46AD] = 8'h00;
RAM[16'h46AE] = 8'h00;
RAM[16'h46AF] = 8'h00;
RAM[16'h46B0] = 8'h00;
RAM[16'h46B1] = 8'h00;
RAM[16'h46B2] = 8'h00;
RAM[16'h46B3] = 8'h00;
RAM[16'h46B4] = 8'h00;
RAM[16'h46B5] = 8'h00;
RAM[16'h46B6] = 8'h00;
RAM[16'h46B7] = 8'h00;
RAM[16'h46B8] = 8'h00;
RAM[16'h46B9] = 8'h00;
RAM[16'h46BA] = 8'h00;
RAM[16'h46BB] = 8'h00;
RAM[16'h46BC] = 8'h00;
RAM[16'h46BD] = 8'h00;
RAM[16'h46BE] = 8'h00;
RAM[16'h46BF] = 8'h00;
RAM[16'h46C0] = 8'h00;
RAM[16'h46C1] = 8'h00;
RAM[16'h46C2] = 8'h00;
RAM[16'h46C3] = 8'h00;
RAM[16'h46C4] = 8'h00;
RAM[16'h46C5] = 8'h00;
RAM[16'h46C6] = 8'h00;
RAM[16'h46C7] = 8'h00;
RAM[16'h46C8] = 8'h00;
RAM[16'h46C9] = 8'h00;
RAM[16'h46CA] = 8'h00;
RAM[16'h46CB] = 8'h00;
RAM[16'h46CC] = 8'h00;
RAM[16'h46CD] = 8'h00;
RAM[16'h46CE] = 8'h00;
RAM[16'h46CF] = 8'h00;
RAM[16'h46D0] = 8'h00;
RAM[16'h46D1] = 8'h00;
RAM[16'h46D2] = 8'h00;
RAM[16'h46D3] = 8'h00;
RAM[16'h46D4] = 8'h00;
RAM[16'h46D5] = 8'h00;
RAM[16'h46D6] = 8'h00;
RAM[16'h46D7] = 8'h00;
RAM[16'h46D8] = 8'h00;
RAM[16'h46D9] = 8'h00;
RAM[16'h46DA] = 8'h00;
RAM[16'h46DB] = 8'h00;
RAM[16'h46DC] = 8'h00;
RAM[16'h46DD] = 8'h00;
RAM[16'h46DE] = 8'h00;
RAM[16'h46DF] = 8'h00;
RAM[16'h46E0] = 8'h00;
RAM[16'h46E1] = 8'h00;
RAM[16'h46E2] = 8'h00;
RAM[16'h46E3] = 8'h00;
RAM[16'h46E4] = 8'h00;
RAM[16'h46E5] = 8'h00;
RAM[16'h46E6] = 8'h00;
RAM[16'h46E7] = 8'h00;
RAM[16'h46E8] = 8'h00;
RAM[16'h46E9] = 8'h00;
RAM[16'h46EA] = 8'h00;
RAM[16'h46EB] = 8'h00;
RAM[16'h46EC] = 8'h00;
RAM[16'h46ED] = 8'h00;
RAM[16'h46EE] = 8'h00;
RAM[16'h46EF] = 8'h00;
RAM[16'h46F0] = 8'h00;
RAM[16'h46F1] = 8'h00;
RAM[16'h46F2] = 8'h00;
RAM[16'h46F3] = 8'h00;
RAM[16'h46F4] = 8'h00;
RAM[16'h46F5] = 8'h00;
RAM[16'h46F6] = 8'h00;
RAM[16'h46F7] = 8'h00;
RAM[16'h46F8] = 8'h00;
RAM[16'h46F9] = 8'h00;
RAM[16'h46FA] = 8'h00;
RAM[16'h46FB] = 8'h00;
RAM[16'h46FC] = 8'h00;
RAM[16'h46FD] = 8'h00;
RAM[16'h46FE] = 8'h00;
RAM[16'h46FF] = 8'h00;
RAM[16'h4700] = 8'h00;
RAM[16'h4701] = 8'h00;
RAM[16'h4702] = 8'h00;
RAM[16'h4703] = 8'h00;
RAM[16'h4704] = 8'h00;
RAM[16'h4705] = 8'h00;
RAM[16'h4706] = 8'h00;
RAM[16'h4707] = 8'h00;
RAM[16'h4708] = 8'h00;
RAM[16'h4709] = 8'h00;
RAM[16'h470A] = 8'h00;
RAM[16'h470B] = 8'h00;
RAM[16'h470C] = 8'h00;
RAM[16'h470D] = 8'h00;
RAM[16'h470E] = 8'h00;
RAM[16'h470F] = 8'h00;
RAM[16'h4710] = 8'h00;
RAM[16'h4711] = 8'h00;
RAM[16'h4712] = 8'h00;
RAM[16'h4713] = 8'h00;
RAM[16'h4714] = 8'h00;
RAM[16'h4715] = 8'h00;
RAM[16'h4716] = 8'h00;
RAM[16'h4717] = 8'h00;
RAM[16'h4718] = 8'h00;
RAM[16'h4719] = 8'h00;
RAM[16'h471A] = 8'h00;
RAM[16'h471B] = 8'h00;
RAM[16'h471C] = 8'h00;
RAM[16'h471D] = 8'h00;
RAM[16'h471E] = 8'h00;
RAM[16'h471F] = 8'h00;
RAM[16'h4720] = 8'h00;
RAM[16'h4721] = 8'h00;
RAM[16'h4722] = 8'h00;
RAM[16'h4723] = 8'h00;
RAM[16'h4724] = 8'h00;
RAM[16'h4725] = 8'h00;
RAM[16'h4726] = 8'h00;
RAM[16'h4727] = 8'h00;
RAM[16'h4728] = 8'h00;
RAM[16'h4729] = 8'h00;
RAM[16'h472A] = 8'h00;
RAM[16'h472B] = 8'h00;
RAM[16'h472C] = 8'h00;
RAM[16'h472D] = 8'h00;
RAM[16'h472E] = 8'h00;
RAM[16'h472F] = 8'h00;
RAM[16'h4730] = 8'h00;
RAM[16'h4731] = 8'h00;
RAM[16'h4732] = 8'h00;
RAM[16'h4733] = 8'h00;
RAM[16'h4734] = 8'h00;
RAM[16'h4735] = 8'h00;
RAM[16'h4736] = 8'h00;
RAM[16'h4737] = 8'h00;
RAM[16'h4738] = 8'h00;
RAM[16'h4739] = 8'h00;
RAM[16'h473A] = 8'h00;
RAM[16'h473B] = 8'h00;
RAM[16'h473C] = 8'h00;
RAM[16'h473D] = 8'h00;
RAM[16'h473E] = 8'h00;
RAM[16'h473F] = 8'h00;
RAM[16'h4740] = 8'h00;
RAM[16'h4741] = 8'h00;
RAM[16'h4742] = 8'h00;
RAM[16'h4743] = 8'h00;
RAM[16'h4744] = 8'h00;
RAM[16'h4745] = 8'h00;
RAM[16'h4746] = 8'h00;
RAM[16'h4747] = 8'h00;
RAM[16'h4748] = 8'h00;
RAM[16'h4749] = 8'h00;
RAM[16'h474A] = 8'h00;
RAM[16'h474B] = 8'h00;
RAM[16'h474C] = 8'h00;
RAM[16'h474D] = 8'h00;
RAM[16'h474E] = 8'h00;
RAM[16'h474F] = 8'h00;
RAM[16'h4750] = 8'h00;
RAM[16'h4751] = 8'h00;
RAM[16'h4752] = 8'h00;
RAM[16'h4753] = 8'h00;
RAM[16'h4754] = 8'h00;
RAM[16'h4755] = 8'h00;
RAM[16'h4756] = 8'h00;
RAM[16'h4757] = 8'h00;
RAM[16'h4758] = 8'h00;
RAM[16'h4759] = 8'h00;
RAM[16'h475A] = 8'h00;
RAM[16'h475B] = 8'h00;
RAM[16'h475C] = 8'h00;
RAM[16'h475D] = 8'h00;
RAM[16'h475E] = 8'h00;
RAM[16'h475F] = 8'h00;
RAM[16'h4760] = 8'h00;
RAM[16'h4761] = 8'h00;
RAM[16'h4762] = 8'h00;
RAM[16'h4763] = 8'h00;
RAM[16'h4764] = 8'h00;
RAM[16'h4765] = 8'h00;
RAM[16'h4766] = 8'h00;
RAM[16'h4767] = 8'h00;
RAM[16'h4768] = 8'h00;
RAM[16'h4769] = 8'h00;
RAM[16'h476A] = 8'h00;
RAM[16'h476B] = 8'h00;
RAM[16'h476C] = 8'h00;
RAM[16'h476D] = 8'h00;
RAM[16'h476E] = 8'h00;
RAM[16'h476F] = 8'h00;
RAM[16'h4770] = 8'h00;
RAM[16'h4771] = 8'h00;
RAM[16'h4772] = 8'h00;
RAM[16'h4773] = 8'h00;
RAM[16'h4774] = 8'h00;
RAM[16'h4775] = 8'h00;
RAM[16'h4776] = 8'h00;
RAM[16'h4777] = 8'h00;
RAM[16'h4778] = 8'h00;
RAM[16'h4779] = 8'h00;
RAM[16'h477A] = 8'h00;
RAM[16'h477B] = 8'h00;
RAM[16'h477C] = 8'h00;
RAM[16'h477D] = 8'h00;
RAM[16'h477E] = 8'h00;
RAM[16'h477F] = 8'h00;
RAM[16'h4780] = 8'h00;
RAM[16'h4781] = 8'h00;
RAM[16'h4782] = 8'h00;
RAM[16'h4783] = 8'h00;
RAM[16'h4784] = 8'h00;
RAM[16'h4785] = 8'h00;
RAM[16'h4786] = 8'h00;
RAM[16'h4787] = 8'h00;
RAM[16'h4788] = 8'h00;
RAM[16'h4789] = 8'h00;
RAM[16'h478A] = 8'h00;
RAM[16'h478B] = 8'h00;
RAM[16'h478C] = 8'h00;
RAM[16'h478D] = 8'h00;
RAM[16'h478E] = 8'h00;
RAM[16'h478F] = 8'h00;
RAM[16'h4790] = 8'h00;
RAM[16'h4791] = 8'h00;
RAM[16'h4792] = 8'h00;
RAM[16'h4793] = 8'h00;
RAM[16'h4794] = 8'h00;
RAM[16'h4795] = 8'h00;
RAM[16'h4796] = 8'h00;
RAM[16'h4797] = 8'h00;
RAM[16'h4798] = 8'h00;
RAM[16'h4799] = 8'h00;
RAM[16'h479A] = 8'h00;
RAM[16'h479B] = 8'h00;
RAM[16'h479C] = 8'h00;
RAM[16'h479D] = 8'h00;
RAM[16'h479E] = 8'h00;
RAM[16'h479F] = 8'h00;
RAM[16'h47A0] = 8'h00;
RAM[16'h47A1] = 8'h00;
RAM[16'h47A2] = 8'h00;
RAM[16'h47A3] = 8'h00;
RAM[16'h47A4] = 8'h00;
RAM[16'h47A5] = 8'h00;
RAM[16'h47A6] = 8'h00;
RAM[16'h47A7] = 8'h00;
RAM[16'h47A8] = 8'h00;
RAM[16'h47A9] = 8'h00;
RAM[16'h47AA] = 8'h00;
RAM[16'h47AB] = 8'h00;
RAM[16'h47AC] = 8'h00;
RAM[16'h47AD] = 8'h00;
RAM[16'h47AE] = 8'h00;
RAM[16'h47AF] = 8'h00;
RAM[16'h47B0] = 8'h00;
RAM[16'h47B1] = 8'h00;
RAM[16'h47B2] = 8'h00;
RAM[16'h47B3] = 8'h00;
RAM[16'h47B4] = 8'h00;
RAM[16'h47B5] = 8'h00;
RAM[16'h47B6] = 8'h00;
RAM[16'h47B7] = 8'h00;
RAM[16'h47B8] = 8'h00;
RAM[16'h47B9] = 8'h00;
RAM[16'h47BA] = 8'h00;
RAM[16'h47BB] = 8'h00;
RAM[16'h47BC] = 8'h00;
RAM[16'h47BD] = 8'h00;
RAM[16'h47BE] = 8'h00;
RAM[16'h47BF] = 8'h00;
RAM[16'h47C0] = 8'h00;
RAM[16'h47C1] = 8'h00;
RAM[16'h47C2] = 8'h00;
RAM[16'h47C3] = 8'h00;
RAM[16'h47C4] = 8'h00;
RAM[16'h47C5] = 8'h00;
RAM[16'h47C6] = 8'h00;
RAM[16'h47C7] = 8'h00;
RAM[16'h47C8] = 8'h00;
RAM[16'h47C9] = 8'h00;
RAM[16'h47CA] = 8'h00;
RAM[16'h47CB] = 8'h00;
RAM[16'h47CC] = 8'h00;
RAM[16'h47CD] = 8'h00;
RAM[16'h47CE] = 8'h00;
RAM[16'h47CF] = 8'h00;
RAM[16'h47D0] = 8'h00;
RAM[16'h47D1] = 8'h00;
RAM[16'h47D2] = 8'h00;
RAM[16'h47D3] = 8'h00;
RAM[16'h47D4] = 8'h00;
RAM[16'h47D5] = 8'h00;
RAM[16'h47D6] = 8'h00;
RAM[16'h47D7] = 8'h00;
RAM[16'h47D8] = 8'h00;
RAM[16'h47D9] = 8'h00;
RAM[16'h47DA] = 8'h00;
RAM[16'h47DB] = 8'h00;
RAM[16'h47DC] = 8'h00;
RAM[16'h47DD] = 8'h00;
RAM[16'h47DE] = 8'h00;
RAM[16'h47DF] = 8'h00;
RAM[16'h47E0] = 8'h00;
RAM[16'h47E1] = 8'h00;
RAM[16'h47E2] = 8'h00;
RAM[16'h47E3] = 8'h00;
RAM[16'h47E4] = 8'h00;
RAM[16'h47E5] = 8'h00;
RAM[16'h47E6] = 8'h00;
RAM[16'h47E7] = 8'h00;
RAM[16'h47E8] = 8'h00;
RAM[16'h47E9] = 8'h00;
RAM[16'h47EA] = 8'h00;
RAM[16'h47EB] = 8'h00;
RAM[16'h47EC] = 8'h00;
RAM[16'h47ED] = 8'h00;
RAM[16'h47EE] = 8'h00;
RAM[16'h47EF] = 8'h00;
RAM[16'h47F0] = 8'h00;
RAM[16'h47F1] = 8'h00;
RAM[16'h47F2] = 8'h00;
RAM[16'h47F3] = 8'h00;
RAM[16'h47F4] = 8'h00;
RAM[16'h47F5] = 8'h00;
RAM[16'h47F6] = 8'h00;
RAM[16'h47F7] = 8'h00;
RAM[16'h47F8] = 8'h00;
RAM[16'h47F9] = 8'h00;
RAM[16'h47FA] = 8'h00;
RAM[16'h47FB] = 8'h00;
RAM[16'h47FC] = 8'h00;
RAM[16'h47FD] = 8'h00;
RAM[16'h47FE] = 8'h00;
RAM[16'h47FF] = 8'h00;
RAM[16'h4800] = 8'h00;
RAM[16'h4801] = 8'h00;
RAM[16'h4802] = 8'h00;
RAM[16'h4803] = 8'h00;
RAM[16'h4804] = 8'h00;
RAM[16'h4805] = 8'h00;
RAM[16'h4806] = 8'h00;
RAM[16'h4807] = 8'h00;
RAM[16'h4808] = 8'h00;
RAM[16'h4809] = 8'h00;
RAM[16'h480A] = 8'h00;
RAM[16'h480B] = 8'h00;
RAM[16'h480C] = 8'h00;
RAM[16'h480D] = 8'h00;
RAM[16'h480E] = 8'h00;
RAM[16'h480F] = 8'h00;
RAM[16'h4810] = 8'h00;
RAM[16'h4811] = 8'h00;
RAM[16'h4812] = 8'h00;
RAM[16'h4813] = 8'h00;
RAM[16'h4814] = 8'h00;
RAM[16'h4815] = 8'h00;
RAM[16'h4816] = 8'h00;
RAM[16'h4817] = 8'h00;
RAM[16'h4818] = 8'h00;
RAM[16'h4819] = 8'h00;
RAM[16'h481A] = 8'h00;
RAM[16'h481B] = 8'h00;
RAM[16'h481C] = 8'h00;
RAM[16'h481D] = 8'h00;
RAM[16'h481E] = 8'h00;
RAM[16'h481F] = 8'h00;
RAM[16'h4820] = 8'h00;
RAM[16'h4821] = 8'h00;
RAM[16'h4822] = 8'h00;
RAM[16'h4823] = 8'h00;
RAM[16'h4824] = 8'h00;
RAM[16'h4825] = 8'h00;
RAM[16'h4826] = 8'h00;
RAM[16'h4827] = 8'h00;
RAM[16'h4828] = 8'h00;
RAM[16'h4829] = 8'h00;
RAM[16'h482A] = 8'h00;
RAM[16'h482B] = 8'h00;
RAM[16'h482C] = 8'h00;
RAM[16'h482D] = 8'h00;
RAM[16'h482E] = 8'h00;
RAM[16'h482F] = 8'h00;
RAM[16'h4830] = 8'h00;
RAM[16'h4831] = 8'h00;
RAM[16'h4832] = 8'h00;
RAM[16'h4833] = 8'h00;
RAM[16'h4834] = 8'h00;
RAM[16'h4835] = 8'h00;
RAM[16'h4836] = 8'h00;
RAM[16'h4837] = 8'h00;
RAM[16'h4838] = 8'h00;
RAM[16'h4839] = 8'h00;
RAM[16'h483A] = 8'h00;
RAM[16'h483B] = 8'h00;
RAM[16'h483C] = 8'h00;
RAM[16'h483D] = 8'h00;
RAM[16'h483E] = 8'h00;
RAM[16'h483F] = 8'h00;
RAM[16'h4840] = 8'h00;
RAM[16'h4841] = 8'h00;
RAM[16'h4842] = 8'h00;
RAM[16'h4843] = 8'h00;
RAM[16'h4844] = 8'h00;
RAM[16'h4845] = 8'h00;
RAM[16'h4846] = 8'h00;
RAM[16'h4847] = 8'h00;
RAM[16'h4848] = 8'h00;
RAM[16'h4849] = 8'h00;
RAM[16'h484A] = 8'h00;
RAM[16'h484B] = 8'h00;
RAM[16'h484C] = 8'h00;
RAM[16'h484D] = 8'h00;
RAM[16'h484E] = 8'h00;
RAM[16'h484F] = 8'h00;
RAM[16'h4850] = 8'h00;
RAM[16'h4851] = 8'h00;
RAM[16'h4852] = 8'h00;
RAM[16'h4853] = 8'h00;
RAM[16'h4854] = 8'h00;
RAM[16'h4855] = 8'h00;
RAM[16'h4856] = 8'h00;
RAM[16'h4857] = 8'h00;
RAM[16'h4858] = 8'h00;
RAM[16'h4859] = 8'h00;
RAM[16'h485A] = 8'h00;
RAM[16'h485B] = 8'h00;
RAM[16'h485C] = 8'h00;
RAM[16'h485D] = 8'h00;
RAM[16'h485E] = 8'h00;
RAM[16'h485F] = 8'h00;
RAM[16'h4860] = 8'h00;
RAM[16'h4861] = 8'h00;
RAM[16'h4862] = 8'h00;
RAM[16'h4863] = 8'h00;
RAM[16'h4864] = 8'h00;
RAM[16'h4865] = 8'h00;
RAM[16'h4866] = 8'h00;
RAM[16'h4867] = 8'h00;
RAM[16'h4868] = 8'h00;
RAM[16'h4869] = 8'h00;
RAM[16'h486A] = 8'h00;
RAM[16'h486B] = 8'h00;
RAM[16'h486C] = 8'h00;
RAM[16'h486D] = 8'h00;
RAM[16'h486E] = 8'h00;
RAM[16'h486F] = 8'h00;
RAM[16'h4870] = 8'h00;
RAM[16'h4871] = 8'h00;
RAM[16'h4872] = 8'h00;
RAM[16'h4873] = 8'h00;
RAM[16'h4874] = 8'h00;
RAM[16'h4875] = 8'h00;
RAM[16'h4876] = 8'h00;
RAM[16'h4877] = 8'h00;
RAM[16'h4878] = 8'h00;
RAM[16'h4879] = 8'h00;
RAM[16'h487A] = 8'h00;
RAM[16'h487B] = 8'h00;
RAM[16'h487C] = 8'h00;
RAM[16'h487D] = 8'h00;
RAM[16'h487E] = 8'h00;
RAM[16'h487F] = 8'h00;
RAM[16'h4880] = 8'h00;
RAM[16'h4881] = 8'h00;
RAM[16'h4882] = 8'h00;
RAM[16'h4883] = 8'h00;
RAM[16'h4884] = 8'h00;
RAM[16'h4885] = 8'h00;
RAM[16'h4886] = 8'h00;
RAM[16'h4887] = 8'h00;
RAM[16'h4888] = 8'h00;
RAM[16'h4889] = 8'h00;
RAM[16'h488A] = 8'h00;
RAM[16'h488B] = 8'h00;
RAM[16'h488C] = 8'h00;
RAM[16'h488D] = 8'h00;
RAM[16'h488E] = 8'h00;
RAM[16'h488F] = 8'h00;
RAM[16'h4890] = 8'h00;
RAM[16'h4891] = 8'h00;
RAM[16'h4892] = 8'h00;
RAM[16'h4893] = 8'h00;
RAM[16'h4894] = 8'h00;
RAM[16'h4895] = 8'h00;
RAM[16'h4896] = 8'h00;
RAM[16'h4897] = 8'h00;
RAM[16'h4898] = 8'h00;
RAM[16'h4899] = 8'h00;
RAM[16'h489A] = 8'h00;
RAM[16'h489B] = 8'h00;
RAM[16'h489C] = 8'h00;
RAM[16'h489D] = 8'h00;
RAM[16'h489E] = 8'h00;
RAM[16'h489F] = 8'h00;
RAM[16'h48A0] = 8'h00;
RAM[16'h48A1] = 8'h00;
RAM[16'h48A2] = 8'h00;
RAM[16'h48A3] = 8'h00;
RAM[16'h48A4] = 8'h00;
RAM[16'h48A5] = 8'h00;
RAM[16'h48A6] = 8'h00;
RAM[16'h48A7] = 8'h00;
RAM[16'h48A8] = 8'h00;
RAM[16'h48A9] = 8'h00;
RAM[16'h48AA] = 8'h00;
RAM[16'h48AB] = 8'h00;
RAM[16'h48AC] = 8'h00;
RAM[16'h48AD] = 8'h00;
RAM[16'h48AE] = 8'h00;
RAM[16'h48AF] = 8'h00;
RAM[16'h48B0] = 8'h00;
RAM[16'h48B1] = 8'h00;
RAM[16'h48B2] = 8'h00;
RAM[16'h48B3] = 8'h00;
RAM[16'h48B4] = 8'h00;
RAM[16'h48B5] = 8'h00;
RAM[16'h48B6] = 8'h00;
RAM[16'h48B7] = 8'h00;
RAM[16'h48B8] = 8'h00;
RAM[16'h48B9] = 8'h00;
RAM[16'h48BA] = 8'h00;
RAM[16'h48BB] = 8'h00;
RAM[16'h48BC] = 8'h00;
RAM[16'h48BD] = 8'h00;
RAM[16'h48BE] = 8'h00;
RAM[16'h48BF] = 8'h00;
RAM[16'h48C0] = 8'h00;
RAM[16'h48C1] = 8'h00;
RAM[16'h48C2] = 8'h00;
RAM[16'h48C3] = 8'h00;
RAM[16'h48C4] = 8'h00;
RAM[16'h48C5] = 8'h00;
RAM[16'h48C6] = 8'h00;
RAM[16'h48C7] = 8'h00;
RAM[16'h48C8] = 8'h00;
RAM[16'h48C9] = 8'h00;
RAM[16'h48CA] = 8'h00;
RAM[16'h48CB] = 8'h00;
RAM[16'h48CC] = 8'h00;
RAM[16'h48CD] = 8'h00;
RAM[16'h48CE] = 8'h00;
RAM[16'h48CF] = 8'h00;
RAM[16'h48D0] = 8'h00;
RAM[16'h48D1] = 8'h00;
RAM[16'h48D2] = 8'h00;
RAM[16'h48D3] = 8'h00;
RAM[16'h48D4] = 8'h00;
RAM[16'h48D5] = 8'h00;
RAM[16'h48D6] = 8'h00;
RAM[16'h48D7] = 8'h00;
RAM[16'h48D8] = 8'h00;
RAM[16'h48D9] = 8'h00;
RAM[16'h48DA] = 8'h00;
RAM[16'h48DB] = 8'h00;
RAM[16'h48DC] = 8'h00;
RAM[16'h48DD] = 8'h00;
RAM[16'h48DE] = 8'h00;
RAM[16'h48DF] = 8'h00;
RAM[16'h48E0] = 8'h00;
RAM[16'h48E1] = 8'h00;
RAM[16'h48E2] = 8'h00;
RAM[16'h48E3] = 8'h00;
RAM[16'h48E4] = 8'h00;
RAM[16'h48E5] = 8'h00;
RAM[16'h48E6] = 8'h00;
RAM[16'h48E7] = 8'h00;
RAM[16'h48E8] = 8'h00;
RAM[16'h48E9] = 8'h00;
RAM[16'h48EA] = 8'h00;
RAM[16'h48EB] = 8'h00;
RAM[16'h48EC] = 8'h00;
RAM[16'h48ED] = 8'h00;
RAM[16'h48EE] = 8'h00;
RAM[16'h48EF] = 8'h00;
RAM[16'h48F0] = 8'h00;
RAM[16'h48F1] = 8'h00;
RAM[16'h48F2] = 8'h00;
RAM[16'h48F3] = 8'h00;
RAM[16'h48F4] = 8'h00;
RAM[16'h48F5] = 8'h00;
RAM[16'h48F6] = 8'h00;
RAM[16'h48F7] = 8'h00;
RAM[16'h48F8] = 8'h00;
RAM[16'h48F9] = 8'h00;
RAM[16'h48FA] = 8'h00;
RAM[16'h48FB] = 8'h00;
RAM[16'h48FC] = 8'h00;
RAM[16'h48FD] = 8'h00;
RAM[16'h48FE] = 8'h00;
RAM[16'h48FF] = 8'h00;
RAM[16'h4900] = 8'h00;
RAM[16'h4901] = 8'h00;
RAM[16'h4902] = 8'h00;
RAM[16'h4903] = 8'h00;
RAM[16'h4904] = 8'h00;
RAM[16'h4905] = 8'h00;
RAM[16'h4906] = 8'h00;
RAM[16'h4907] = 8'h00;
RAM[16'h4908] = 8'h00;
RAM[16'h4909] = 8'h00;
RAM[16'h490A] = 8'h00;
RAM[16'h490B] = 8'h00;
RAM[16'h490C] = 8'h00;
RAM[16'h490D] = 8'h00;
RAM[16'h490E] = 8'h00;
RAM[16'h490F] = 8'h00;
RAM[16'h4910] = 8'h00;
RAM[16'h4911] = 8'h00;
RAM[16'h4912] = 8'h00;
RAM[16'h4913] = 8'h00;
RAM[16'h4914] = 8'h00;
RAM[16'h4915] = 8'h00;
RAM[16'h4916] = 8'h00;
RAM[16'h4917] = 8'h00;
RAM[16'h4918] = 8'h00;
RAM[16'h4919] = 8'h00;
RAM[16'h491A] = 8'h00;
RAM[16'h491B] = 8'h00;
RAM[16'h491C] = 8'h00;
RAM[16'h491D] = 8'h00;
RAM[16'h491E] = 8'h00;
RAM[16'h491F] = 8'h00;
RAM[16'h4920] = 8'h00;
RAM[16'h4921] = 8'h00;
RAM[16'h4922] = 8'h00;
RAM[16'h4923] = 8'h00;
RAM[16'h4924] = 8'h00;
RAM[16'h4925] = 8'h00;
RAM[16'h4926] = 8'h00;
RAM[16'h4927] = 8'h00;
RAM[16'h4928] = 8'h00;
RAM[16'h4929] = 8'h00;
RAM[16'h492A] = 8'h00;
RAM[16'h492B] = 8'h00;
RAM[16'h492C] = 8'h00;
RAM[16'h492D] = 8'h00;
RAM[16'h492E] = 8'h00;
RAM[16'h492F] = 8'h00;
RAM[16'h4930] = 8'h00;
RAM[16'h4931] = 8'h00;
RAM[16'h4932] = 8'h00;
RAM[16'h4933] = 8'h00;
RAM[16'h4934] = 8'h00;
RAM[16'h4935] = 8'h00;
RAM[16'h4936] = 8'h00;
RAM[16'h4937] = 8'h00;
RAM[16'h4938] = 8'h00;
RAM[16'h4939] = 8'h00;
RAM[16'h493A] = 8'h00;
RAM[16'h493B] = 8'h00;
RAM[16'h493C] = 8'h00;
RAM[16'h493D] = 8'h00;
RAM[16'h493E] = 8'h00;
RAM[16'h493F] = 8'h00;
RAM[16'h4940] = 8'h00;
RAM[16'h4941] = 8'h00;
RAM[16'h4942] = 8'h00;
RAM[16'h4943] = 8'h00;
RAM[16'h4944] = 8'h00;
RAM[16'h4945] = 8'h00;
RAM[16'h4946] = 8'h00;
RAM[16'h4947] = 8'h00;
RAM[16'h4948] = 8'h00;
RAM[16'h4949] = 8'h00;
RAM[16'h494A] = 8'h00;
RAM[16'h494B] = 8'h00;
RAM[16'h494C] = 8'h00;
RAM[16'h494D] = 8'h00;
RAM[16'h494E] = 8'h00;
RAM[16'h494F] = 8'h00;
RAM[16'h4950] = 8'h00;
RAM[16'h4951] = 8'h00;
RAM[16'h4952] = 8'h00;
RAM[16'h4953] = 8'h00;
RAM[16'h4954] = 8'h00;
RAM[16'h4955] = 8'h00;
RAM[16'h4956] = 8'h00;
RAM[16'h4957] = 8'h00;
RAM[16'h4958] = 8'h00;
RAM[16'h4959] = 8'h00;
RAM[16'h495A] = 8'h00;
RAM[16'h495B] = 8'h00;
RAM[16'h495C] = 8'h00;
RAM[16'h495D] = 8'h00;
RAM[16'h495E] = 8'h00;
RAM[16'h495F] = 8'h00;
RAM[16'h4960] = 8'h00;
RAM[16'h4961] = 8'h00;
RAM[16'h4962] = 8'h00;
RAM[16'h4963] = 8'h00;
RAM[16'h4964] = 8'h00;
RAM[16'h4965] = 8'h00;
RAM[16'h4966] = 8'h00;
RAM[16'h4967] = 8'h00;
RAM[16'h4968] = 8'h00;
RAM[16'h4969] = 8'h00;
RAM[16'h496A] = 8'h00;
RAM[16'h496B] = 8'h00;
RAM[16'h496C] = 8'h00;
RAM[16'h496D] = 8'h00;
RAM[16'h496E] = 8'h00;
RAM[16'h496F] = 8'h00;
RAM[16'h4970] = 8'h00;
RAM[16'h4971] = 8'h00;
RAM[16'h4972] = 8'h00;
RAM[16'h4973] = 8'h00;
RAM[16'h4974] = 8'h00;
RAM[16'h4975] = 8'h00;
RAM[16'h4976] = 8'h00;
RAM[16'h4977] = 8'h00;
RAM[16'h4978] = 8'h00;
RAM[16'h4979] = 8'h00;
RAM[16'h497A] = 8'h00;
RAM[16'h497B] = 8'h00;
RAM[16'h497C] = 8'h00;
RAM[16'h497D] = 8'h00;
RAM[16'h497E] = 8'h00;
RAM[16'h497F] = 8'h00;
RAM[16'h4980] = 8'h00;
RAM[16'h4981] = 8'h00;
RAM[16'h4982] = 8'h00;
RAM[16'h4983] = 8'h00;
RAM[16'h4984] = 8'h00;
RAM[16'h4985] = 8'h00;
RAM[16'h4986] = 8'h00;
RAM[16'h4987] = 8'h00;
RAM[16'h4988] = 8'h00;
RAM[16'h4989] = 8'h00;
RAM[16'h498A] = 8'h00;
RAM[16'h498B] = 8'h00;
RAM[16'h498C] = 8'h00;
RAM[16'h498D] = 8'h00;
RAM[16'h498E] = 8'h00;
RAM[16'h498F] = 8'h00;
RAM[16'h4990] = 8'h00;
RAM[16'h4991] = 8'h00;
RAM[16'h4992] = 8'h00;
RAM[16'h4993] = 8'h00;
RAM[16'h4994] = 8'h00;
RAM[16'h4995] = 8'h00;
RAM[16'h4996] = 8'h00;
RAM[16'h4997] = 8'h00;
RAM[16'h4998] = 8'h00;
RAM[16'h4999] = 8'h00;
RAM[16'h499A] = 8'h00;
RAM[16'h499B] = 8'h00;
RAM[16'h499C] = 8'h00;
RAM[16'h499D] = 8'h00;
RAM[16'h499E] = 8'h00;
RAM[16'h499F] = 8'h00;
RAM[16'h49A0] = 8'h00;
RAM[16'h49A1] = 8'h00;
RAM[16'h49A2] = 8'h00;
RAM[16'h49A3] = 8'h00;
RAM[16'h49A4] = 8'h00;
RAM[16'h49A5] = 8'h00;
RAM[16'h49A6] = 8'h00;
RAM[16'h49A7] = 8'h00;
RAM[16'h49A8] = 8'h00;
RAM[16'h49A9] = 8'h00;
RAM[16'h49AA] = 8'h00;
RAM[16'h49AB] = 8'h00;
RAM[16'h49AC] = 8'h00;
RAM[16'h49AD] = 8'h00;
RAM[16'h49AE] = 8'h00;
RAM[16'h49AF] = 8'h00;
RAM[16'h49B0] = 8'h00;
RAM[16'h49B1] = 8'h00;
RAM[16'h49B2] = 8'h00;
RAM[16'h49B3] = 8'h00;
RAM[16'h49B4] = 8'h00;
RAM[16'h49B5] = 8'h00;
RAM[16'h49B6] = 8'h00;
RAM[16'h49B7] = 8'h00;
RAM[16'h49B8] = 8'h00;
RAM[16'h49B9] = 8'h00;
RAM[16'h49BA] = 8'h00;
RAM[16'h49BB] = 8'h00;
RAM[16'h49BC] = 8'h00;
RAM[16'h49BD] = 8'h00;
RAM[16'h49BE] = 8'h00;
RAM[16'h49BF] = 8'h00;
RAM[16'h49C0] = 8'h00;
RAM[16'h49C1] = 8'h00;
RAM[16'h49C2] = 8'h00;
RAM[16'h49C3] = 8'h00;
RAM[16'h49C4] = 8'h00;
RAM[16'h49C5] = 8'h00;
RAM[16'h49C6] = 8'h00;
RAM[16'h49C7] = 8'h00;
RAM[16'h49C8] = 8'h00;
RAM[16'h49C9] = 8'h00;
RAM[16'h49CA] = 8'h00;
RAM[16'h49CB] = 8'h00;
RAM[16'h49CC] = 8'h00;
RAM[16'h49CD] = 8'h00;
RAM[16'h49CE] = 8'h00;
RAM[16'h49CF] = 8'h00;
RAM[16'h49D0] = 8'h00;
RAM[16'h49D1] = 8'h00;
RAM[16'h49D2] = 8'h00;
RAM[16'h49D3] = 8'h00;
RAM[16'h49D4] = 8'h00;
RAM[16'h49D5] = 8'h00;
RAM[16'h49D6] = 8'h00;
RAM[16'h49D7] = 8'h00;
RAM[16'h49D8] = 8'h00;
RAM[16'h49D9] = 8'h00;
RAM[16'h49DA] = 8'h00;
RAM[16'h49DB] = 8'h00;
RAM[16'h49DC] = 8'h00;
RAM[16'h49DD] = 8'h00;
RAM[16'h49DE] = 8'h00;
RAM[16'h49DF] = 8'h00;
RAM[16'h49E0] = 8'h00;
RAM[16'h49E1] = 8'h00;
RAM[16'h49E2] = 8'h00;
RAM[16'h49E3] = 8'h00;
RAM[16'h49E4] = 8'h00;
RAM[16'h49E5] = 8'h00;
RAM[16'h49E6] = 8'h00;
RAM[16'h49E7] = 8'h00;
RAM[16'h49E8] = 8'h00;
RAM[16'h49E9] = 8'h00;
RAM[16'h49EA] = 8'h00;
RAM[16'h49EB] = 8'h00;
RAM[16'h49EC] = 8'h00;
RAM[16'h49ED] = 8'h00;
RAM[16'h49EE] = 8'h00;
RAM[16'h49EF] = 8'h00;
RAM[16'h49F0] = 8'h00;
RAM[16'h49F1] = 8'h00;
RAM[16'h49F2] = 8'h00;
RAM[16'h49F3] = 8'h00;
RAM[16'h49F4] = 8'h00;
RAM[16'h49F5] = 8'h00;
RAM[16'h49F6] = 8'h00;
RAM[16'h49F7] = 8'h00;
RAM[16'h49F8] = 8'h00;
RAM[16'h49F9] = 8'h00;
RAM[16'h49FA] = 8'h00;
RAM[16'h49FB] = 8'h00;
RAM[16'h49FC] = 8'h00;
RAM[16'h49FD] = 8'h00;
RAM[16'h49FE] = 8'h00;
RAM[16'h49FF] = 8'h00;
RAM[16'h4A00] = 8'h00;
RAM[16'h4A01] = 8'h00;
RAM[16'h4A02] = 8'h00;
RAM[16'h4A03] = 8'h00;
RAM[16'h4A04] = 8'h00;
RAM[16'h4A05] = 8'h00;
RAM[16'h4A06] = 8'h00;
RAM[16'h4A07] = 8'h00;
RAM[16'h4A08] = 8'h00;
RAM[16'h4A09] = 8'h00;
RAM[16'h4A0A] = 8'h00;
RAM[16'h4A0B] = 8'h00;
RAM[16'h4A0C] = 8'h00;
RAM[16'h4A0D] = 8'h00;
RAM[16'h4A0E] = 8'h00;
RAM[16'h4A0F] = 8'h00;
RAM[16'h4A10] = 8'h00;
RAM[16'h4A11] = 8'h00;
RAM[16'h4A12] = 8'h00;
RAM[16'h4A13] = 8'h00;
RAM[16'h4A14] = 8'h00;
RAM[16'h4A15] = 8'h00;
RAM[16'h4A16] = 8'h00;
RAM[16'h4A17] = 8'h00;
RAM[16'h4A18] = 8'h00;
RAM[16'h4A19] = 8'h00;
RAM[16'h4A1A] = 8'h00;
RAM[16'h4A1B] = 8'h00;
RAM[16'h4A1C] = 8'h00;
RAM[16'h4A1D] = 8'h00;
RAM[16'h4A1E] = 8'h00;
RAM[16'h4A1F] = 8'h00;
RAM[16'h4A20] = 8'h00;
RAM[16'h4A21] = 8'h00;
RAM[16'h4A22] = 8'h00;
RAM[16'h4A23] = 8'h00;
RAM[16'h4A24] = 8'h00;
RAM[16'h4A25] = 8'h00;
RAM[16'h4A26] = 8'h00;
RAM[16'h4A27] = 8'h00;
RAM[16'h4A28] = 8'h00;
RAM[16'h4A29] = 8'h00;
RAM[16'h4A2A] = 8'h00;
RAM[16'h4A2B] = 8'h00;
RAM[16'h4A2C] = 8'h00;
RAM[16'h4A2D] = 8'h00;
RAM[16'h4A2E] = 8'h00;
RAM[16'h4A2F] = 8'h00;
RAM[16'h4A30] = 8'h00;
RAM[16'h4A31] = 8'h00;
RAM[16'h4A32] = 8'h00;
RAM[16'h4A33] = 8'h00;
RAM[16'h4A34] = 8'h00;
RAM[16'h4A35] = 8'h00;
RAM[16'h4A36] = 8'h00;
RAM[16'h4A37] = 8'h00;
RAM[16'h4A38] = 8'h00;
RAM[16'h4A39] = 8'h00;
RAM[16'h4A3A] = 8'h00;
RAM[16'h4A3B] = 8'h00;
RAM[16'h4A3C] = 8'h00;
RAM[16'h4A3D] = 8'h00;
RAM[16'h4A3E] = 8'h00;
RAM[16'h4A3F] = 8'h00;
RAM[16'h4A40] = 8'h00;
RAM[16'h4A41] = 8'h00;
RAM[16'h4A42] = 8'h00;
RAM[16'h4A43] = 8'h00;
RAM[16'h4A44] = 8'h00;
RAM[16'h4A45] = 8'h00;
RAM[16'h4A46] = 8'h00;
RAM[16'h4A47] = 8'h00;
RAM[16'h4A48] = 8'h00;
RAM[16'h4A49] = 8'h00;
RAM[16'h4A4A] = 8'h00;
RAM[16'h4A4B] = 8'h00;
RAM[16'h4A4C] = 8'h00;
RAM[16'h4A4D] = 8'h00;
RAM[16'h4A4E] = 8'h00;
RAM[16'h4A4F] = 8'h00;
RAM[16'h4A50] = 8'h00;
RAM[16'h4A51] = 8'h00;
RAM[16'h4A52] = 8'h00;
RAM[16'h4A53] = 8'h00;
RAM[16'h4A54] = 8'h00;
RAM[16'h4A55] = 8'h00;
RAM[16'h4A56] = 8'h00;
RAM[16'h4A57] = 8'h00;
RAM[16'h4A58] = 8'h00;
RAM[16'h4A59] = 8'h00;
RAM[16'h4A5A] = 8'h00;
RAM[16'h4A5B] = 8'h00;
RAM[16'h4A5C] = 8'h00;
RAM[16'h4A5D] = 8'h00;
RAM[16'h4A5E] = 8'h00;
RAM[16'h4A5F] = 8'h00;
RAM[16'h4A60] = 8'h00;
RAM[16'h4A61] = 8'h00;
RAM[16'h4A62] = 8'h00;
RAM[16'h4A63] = 8'h00;
RAM[16'h4A64] = 8'h00;
RAM[16'h4A65] = 8'h00;
RAM[16'h4A66] = 8'h00;
RAM[16'h4A67] = 8'h00;
RAM[16'h4A68] = 8'h00;
RAM[16'h4A69] = 8'h00;
RAM[16'h4A6A] = 8'h00;
RAM[16'h4A6B] = 8'h00;
RAM[16'h4A6C] = 8'h00;
RAM[16'h4A6D] = 8'h00;
RAM[16'h4A6E] = 8'h00;
RAM[16'h4A6F] = 8'h00;
RAM[16'h4A70] = 8'h00;
RAM[16'h4A71] = 8'h00;
RAM[16'h4A72] = 8'h00;
RAM[16'h4A73] = 8'h00;
RAM[16'h4A74] = 8'h00;
RAM[16'h4A75] = 8'h00;
RAM[16'h4A76] = 8'h00;
RAM[16'h4A77] = 8'h00;
RAM[16'h4A78] = 8'h00;
RAM[16'h4A79] = 8'h00;
RAM[16'h4A7A] = 8'h00;
RAM[16'h4A7B] = 8'h00;
RAM[16'h4A7C] = 8'h00;
RAM[16'h4A7D] = 8'h00;
RAM[16'h4A7E] = 8'h00;
RAM[16'h4A7F] = 8'h00;
RAM[16'h4A80] = 8'h00;
RAM[16'h4A81] = 8'h00;
RAM[16'h4A82] = 8'h00;
RAM[16'h4A83] = 8'h00;
RAM[16'h4A84] = 8'h00;
RAM[16'h4A85] = 8'h00;
RAM[16'h4A86] = 8'h00;
RAM[16'h4A87] = 8'h00;
RAM[16'h4A88] = 8'h00;
RAM[16'h4A89] = 8'h00;
RAM[16'h4A8A] = 8'h00;
RAM[16'h4A8B] = 8'h00;
RAM[16'h4A8C] = 8'h00;
RAM[16'h4A8D] = 8'h00;
RAM[16'h4A8E] = 8'h00;
RAM[16'h4A8F] = 8'h00;
RAM[16'h4A90] = 8'h00;
RAM[16'h4A91] = 8'h00;
RAM[16'h4A92] = 8'h00;
RAM[16'h4A93] = 8'h00;
RAM[16'h4A94] = 8'h00;
RAM[16'h4A95] = 8'h00;
RAM[16'h4A96] = 8'h00;
RAM[16'h4A97] = 8'h00;
RAM[16'h4A98] = 8'h00;
RAM[16'h4A99] = 8'h00;
RAM[16'h4A9A] = 8'h00;
RAM[16'h4A9B] = 8'h00;
RAM[16'h4A9C] = 8'h00;
RAM[16'h4A9D] = 8'h00;
RAM[16'h4A9E] = 8'h00;
RAM[16'h4A9F] = 8'h00;
RAM[16'h4AA0] = 8'h00;
RAM[16'h4AA1] = 8'h00;
RAM[16'h4AA2] = 8'h00;
RAM[16'h4AA3] = 8'h00;
RAM[16'h4AA4] = 8'h00;
RAM[16'h4AA5] = 8'h00;
RAM[16'h4AA6] = 8'h00;
RAM[16'h4AA7] = 8'h00;
RAM[16'h4AA8] = 8'h00;
RAM[16'h4AA9] = 8'h00;
RAM[16'h4AAA] = 8'h00;
RAM[16'h4AAB] = 8'h00;
RAM[16'h4AAC] = 8'h00;
RAM[16'h4AAD] = 8'h00;
RAM[16'h4AAE] = 8'h00;
RAM[16'h4AAF] = 8'h00;
RAM[16'h4AB0] = 8'h00;
RAM[16'h4AB1] = 8'h00;
RAM[16'h4AB2] = 8'h00;
RAM[16'h4AB3] = 8'h00;
RAM[16'h4AB4] = 8'h00;
RAM[16'h4AB5] = 8'h00;
RAM[16'h4AB6] = 8'h00;
RAM[16'h4AB7] = 8'h00;
RAM[16'h4AB8] = 8'h00;
RAM[16'h4AB9] = 8'h00;
RAM[16'h4ABA] = 8'h00;
RAM[16'h4ABB] = 8'h00;
RAM[16'h4ABC] = 8'h00;
RAM[16'h4ABD] = 8'h00;
RAM[16'h4ABE] = 8'h00;
RAM[16'h4ABF] = 8'h00;
RAM[16'h4AC0] = 8'h00;
RAM[16'h4AC1] = 8'h00;
RAM[16'h4AC2] = 8'h00;
RAM[16'h4AC3] = 8'h00;
RAM[16'h4AC4] = 8'h00;
RAM[16'h4AC5] = 8'h00;
RAM[16'h4AC6] = 8'h00;
RAM[16'h4AC7] = 8'h00;
RAM[16'h4AC8] = 8'h00;
RAM[16'h4AC9] = 8'h00;
RAM[16'h4ACA] = 8'h00;
RAM[16'h4ACB] = 8'h00;
RAM[16'h4ACC] = 8'h00;
RAM[16'h4ACD] = 8'h00;
RAM[16'h4ACE] = 8'h00;
RAM[16'h4ACF] = 8'h00;
RAM[16'h4AD0] = 8'h00;
RAM[16'h4AD1] = 8'h00;
RAM[16'h4AD2] = 8'h00;
RAM[16'h4AD3] = 8'h00;
RAM[16'h4AD4] = 8'h00;
RAM[16'h4AD5] = 8'h00;
RAM[16'h4AD6] = 8'h00;
RAM[16'h4AD7] = 8'h00;
RAM[16'h4AD8] = 8'h00;
RAM[16'h4AD9] = 8'h00;
RAM[16'h4ADA] = 8'h00;
RAM[16'h4ADB] = 8'h00;
RAM[16'h4ADC] = 8'h00;
RAM[16'h4ADD] = 8'h00;
RAM[16'h4ADE] = 8'h00;
RAM[16'h4ADF] = 8'h00;
RAM[16'h4AE0] = 8'h00;
RAM[16'h4AE1] = 8'h00;
RAM[16'h4AE2] = 8'h00;
RAM[16'h4AE3] = 8'h00;
RAM[16'h4AE4] = 8'h00;
RAM[16'h4AE5] = 8'h00;
RAM[16'h4AE6] = 8'h00;
RAM[16'h4AE7] = 8'h00;
RAM[16'h4AE8] = 8'h00;
RAM[16'h4AE9] = 8'h00;
RAM[16'h4AEA] = 8'h00;
RAM[16'h4AEB] = 8'h00;
RAM[16'h4AEC] = 8'h00;
RAM[16'h4AED] = 8'h00;
RAM[16'h4AEE] = 8'h00;
RAM[16'h4AEF] = 8'h00;
RAM[16'h4AF0] = 8'h00;
RAM[16'h4AF1] = 8'h00;
RAM[16'h4AF2] = 8'h00;
RAM[16'h4AF3] = 8'h00;
RAM[16'h4AF4] = 8'h00;
RAM[16'h4AF5] = 8'h00;
RAM[16'h4AF6] = 8'h00;
RAM[16'h4AF7] = 8'h00;
RAM[16'h4AF8] = 8'h00;
RAM[16'h4AF9] = 8'h00;
RAM[16'h4AFA] = 8'h00;
RAM[16'h4AFB] = 8'h00;
RAM[16'h4AFC] = 8'h00;
RAM[16'h4AFD] = 8'h00;
RAM[16'h4AFE] = 8'h00;
RAM[16'h4AFF] = 8'h00;
RAM[16'h4B00] = 8'h00;
RAM[16'h4B01] = 8'h00;
RAM[16'h4B02] = 8'h00;
RAM[16'h4B03] = 8'h00;
RAM[16'h4B04] = 8'h00;
RAM[16'h4B05] = 8'h00;
RAM[16'h4B06] = 8'h00;
RAM[16'h4B07] = 8'h00;
RAM[16'h4B08] = 8'h00;
RAM[16'h4B09] = 8'h00;
RAM[16'h4B0A] = 8'h00;
RAM[16'h4B0B] = 8'h00;
RAM[16'h4B0C] = 8'h00;
RAM[16'h4B0D] = 8'h00;
RAM[16'h4B0E] = 8'h00;
RAM[16'h4B0F] = 8'h00;
RAM[16'h4B10] = 8'h00;
RAM[16'h4B11] = 8'h00;
RAM[16'h4B12] = 8'h00;
RAM[16'h4B13] = 8'h00;
RAM[16'h4B14] = 8'h00;
RAM[16'h4B15] = 8'h00;
RAM[16'h4B16] = 8'h00;
RAM[16'h4B17] = 8'h00;
RAM[16'h4B18] = 8'h00;
RAM[16'h4B19] = 8'h00;
RAM[16'h4B1A] = 8'h00;
RAM[16'h4B1B] = 8'h00;
RAM[16'h4B1C] = 8'h00;
RAM[16'h4B1D] = 8'h00;
RAM[16'h4B1E] = 8'h00;
RAM[16'h4B1F] = 8'h00;
RAM[16'h4B20] = 8'h00;
RAM[16'h4B21] = 8'h00;
RAM[16'h4B22] = 8'h00;
RAM[16'h4B23] = 8'h00;
RAM[16'h4B24] = 8'h00;
RAM[16'h4B25] = 8'h00;
RAM[16'h4B26] = 8'h00;
RAM[16'h4B27] = 8'h00;
RAM[16'h4B28] = 8'h00;
RAM[16'h4B29] = 8'h00;
RAM[16'h4B2A] = 8'h00;
RAM[16'h4B2B] = 8'h00;
RAM[16'h4B2C] = 8'h00;
RAM[16'h4B2D] = 8'h00;
RAM[16'h4B2E] = 8'h00;
RAM[16'h4B2F] = 8'h00;
RAM[16'h4B30] = 8'h00;
RAM[16'h4B31] = 8'h00;
RAM[16'h4B32] = 8'h00;
RAM[16'h4B33] = 8'h00;
RAM[16'h4B34] = 8'h00;
RAM[16'h4B35] = 8'h00;
RAM[16'h4B36] = 8'h00;
RAM[16'h4B37] = 8'h00;
RAM[16'h4B38] = 8'h00;
RAM[16'h4B39] = 8'h00;
RAM[16'h4B3A] = 8'h00;
RAM[16'h4B3B] = 8'h00;
RAM[16'h4B3C] = 8'h00;
RAM[16'h4B3D] = 8'h00;
RAM[16'h4B3E] = 8'h00;
RAM[16'h4B3F] = 8'h00;
RAM[16'h4B40] = 8'h00;
RAM[16'h4B41] = 8'h00;
RAM[16'h4B42] = 8'h00;
RAM[16'h4B43] = 8'h00;
RAM[16'h4B44] = 8'h00;
RAM[16'h4B45] = 8'h00;
RAM[16'h4B46] = 8'h00;
RAM[16'h4B47] = 8'h00;
RAM[16'h4B48] = 8'h00;
RAM[16'h4B49] = 8'h00;
RAM[16'h4B4A] = 8'h00;
RAM[16'h4B4B] = 8'h00;
RAM[16'h4B4C] = 8'h00;
RAM[16'h4B4D] = 8'h00;
RAM[16'h4B4E] = 8'h00;
RAM[16'h4B4F] = 8'h00;
RAM[16'h4B50] = 8'h00;
RAM[16'h4B51] = 8'h00;
RAM[16'h4B52] = 8'h00;
RAM[16'h4B53] = 8'h00;
RAM[16'h4B54] = 8'h00;
RAM[16'h4B55] = 8'h00;
RAM[16'h4B56] = 8'h00;
RAM[16'h4B57] = 8'h00;
RAM[16'h4B58] = 8'h00;
RAM[16'h4B59] = 8'h00;
RAM[16'h4B5A] = 8'h00;
RAM[16'h4B5B] = 8'h00;
RAM[16'h4B5C] = 8'h00;
RAM[16'h4B5D] = 8'h00;
RAM[16'h4B5E] = 8'h00;
RAM[16'h4B5F] = 8'h00;
RAM[16'h4B60] = 8'h00;
RAM[16'h4B61] = 8'h00;
RAM[16'h4B62] = 8'h00;
RAM[16'h4B63] = 8'h00;
RAM[16'h4B64] = 8'h00;
RAM[16'h4B65] = 8'h00;
RAM[16'h4B66] = 8'h00;
RAM[16'h4B67] = 8'h00;
RAM[16'h4B68] = 8'h00;
RAM[16'h4B69] = 8'h00;
RAM[16'h4B6A] = 8'h00;
RAM[16'h4B6B] = 8'h00;
RAM[16'h4B6C] = 8'h00;
RAM[16'h4B6D] = 8'h00;
RAM[16'h4B6E] = 8'h00;
RAM[16'h4B6F] = 8'h00;
RAM[16'h4B70] = 8'h00;
RAM[16'h4B71] = 8'h00;
RAM[16'h4B72] = 8'h00;
RAM[16'h4B73] = 8'h00;
RAM[16'h4B74] = 8'h00;
RAM[16'h4B75] = 8'h00;
RAM[16'h4B76] = 8'h00;
RAM[16'h4B77] = 8'h00;
RAM[16'h4B78] = 8'h00;
RAM[16'h4B79] = 8'h00;
RAM[16'h4B7A] = 8'h00;
RAM[16'h4B7B] = 8'h00;
RAM[16'h4B7C] = 8'h00;
RAM[16'h4B7D] = 8'h00;
RAM[16'h4B7E] = 8'h00;
RAM[16'h4B7F] = 8'h00;
RAM[16'h4B80] = 8'h00;
RAM[16'h4B81] = 8'h00;
RAM[16'h4B82] = 8'h00;
RAM[16'h4B83] = 8'h00;
RAM[16'h4B84] = 8'h00;
RAM[16'h4B85] = 8'h00;
RAM[16'h4B86] = 8'h00;
RAM[16'h4B87] = 8'h00;
RAM[16'h4B88] = 8'h00;
RAM[16'h4B89] = 8'h00;
RAM[16'h4B8A] = 8'h00;
RAM[16'h4B8B] = 8'h00;
RAM[16'h4B8C] = 8'h00;
RAM[16'h4B8D] = 8'h00;
RAM[16'h4B8E] = 8'h00;
RAM[16'h4B8F] = 8'h00;
RAM[16'h4B90] = 8'h00;
RAM[16'h4B91] = 8'h00;
RAM[16'h4B92] = 8'h00;
RAM[16'h4B93] = 8'h00;
RAM[16'h4B94] = 8'h00;
RAM[16'h4B95] = 8'h00;
RAM[16'h4B96] = 8'h00;
RAM[16'h4B97] = 8'h00;
RAM[16'h4B98] = 8'h00;
RAM[16'h4B99] = 8'h00;
RAM[16'h4B9A] = 8'h00;
RAM[16'h4B9B] = 8'h00;
RAM[16'h4B9C] = 8'h00;
RAM[16'h4B9D] = 8'h00;
RAM[16'h4B9E] = 8'h00;
RAM[16'h4B9F] = 8'h00;
RAM[16'h4BA0] = 8'h00;
RAM[16'h4BA1] = 8'h00;
RAM[16'h4BA2] = 8'h00;
RAM[16'h4BA3] = 8'h00;
RAM[16'h4BA4] = 8'h00;
RAM[16'h4BA5] = 8'h00;
RAM[16'h4BA6] = 8'h00;
RAM[16'h4BA7] = 8'h00;
RAM[16'h4BA8] = 8'h00;
RAM[16'h4BA9] = 8'h00;
RAM[16'h4BAA] = 8'h00;
RAM[16'h4BAB] = 8'h00;
RAM[16'h4BAC] = 8'h00;
RAM[16'h4BAD] = 8'h00;
RAM[16'h4BAE] = 8'h00;
RAM[16'h4BAF] = 8'h00;
RAM[16'h4BB0] = 8'h00;
RAM[16'h4BB1] = 8'h00;
RAM[16'h4BB2] = 8'h00;
RAM[16'h4BB3] = 8'h00;
RAM[16'h4BB4] = 8'h00;
RAM[16'h4BB5] = 8'h00;
RAM[16'h4BB6] = 8'h00;
RAM[16'h4BB7] = 8'h00;
RAM[16'h4BB8] = 8'h00;
RAM[16'h4BB9] = 8'h00;
RAM[16'h4BBA] = 8'h00;
RAM[16'h4BBB] = 8'h00;
RAM[16'h4BBC] = 8'h00;
RAM[16'h4BBD] = 8'h00;
RAM[16'h4BBE] = 8'h00;
RAM[16'h4BBF] = 8'h00;
RAM[16'h4BC0] = 8'h00;
RAM[16'h4BC1] = 8'h00;
RAM[16'h4BC2] = 8'h00;
RAM[16'h4BC3] = 8'h00;
RAM[16'h4BC4] = 8'h00;
RAM[16'h4BC5] = 8'h00;
RAM[16'h4BC6] = 8'h00;
RAM[16'h4BC7] = 8'h00;
RAM[16'h4BC8] = 8'h00;
RAM[16'h4BC9] = 8'h00;
RAM[16'h4BCA] = 8'h00;
RAM[16'h4BCB] = 8'h00;
RAM[16'h4BCC] = 8'h00;
RAM[16'h4BCD] = 8'h00;
RAM[16'h4BCE] = 8'h00;
RAM[16'h4BCF] = 8'h00;
RAM[16'h4BD0] = 8'h00;
RAM[16'h4BD1] = 8'h00;
RAM[16'h4BD2] = 8'h00;
RAM[16'h4BD3] = 8'h00;
RAM[16'h4BD4] = 8'h00;
RAM[16'h4BD5] = 8'h00;
RAM[16'h4BD6] = 8'h00;
RAM[16'h4BD7] = 8'h00;
RAM[16'h4BD8] = 8'h00;
RAM[16'h4BD9] = 8'h00;
RAM[16'h4BDA] = 8'h00;
RAM[16'h4BDB] = 8'h00;
RAM[16'h4BDC] = 8'h00;
RAM[16'h4BDD] = 8'h00;
RAM[16'h4BDE] = 8'h00;
RAM[16'h4BDF] = 8'h00;
RAM[16'h4BE0] = 8'h00;
RAM[16'h4BE1] = 8'h00;
RAM[16'h4BE2] = 8'h00;
RAM[16'h4BE3] = 8'h00;
RAM[16'h4BE4] = 8'h00;
RAM[16'h4BE5] = 8'h00;
RAM[16'h4BE6] = 8'h00;
RAM[16'h4BE7] = 8'h00;
RAM[16'h4BE8] = 8'h00;
RAM[16'h4BE9] = 8'h00;
RAM[16'h4BEA] = 8'h00;
RAM[16'h4BEB] = 8'h00;
RAM[16'h4BEC] = 8'h00;
RAM[16'h4BED] = 8'h00;
RAM[16'h4BEE] = 8'h00;
RAM[16'h4BEF] = 8'h00;
RAM[16'h4BF0] = 8'h00;
RAM[16'h4BF1] = 8'h00;
RAM[16'h4BF2] = 8'h00;
RAM[16'h4BF3] = 8'h00;
RAM[16'h4BF4] = 8'h00;
RAM[16'h4BF5] = 8'h00;
RAM[16'h4BF6] = 8'h00;
RAM[16'h4BF7] = 8'h00;
RAM[16'h4BF8] = 8'h00;
RAM[16'h4BF9] = 8'h00;
RAM[16'h4BFA] = 8'h00;
RAM[16'h4BFB] = 8'h00;
RAM[16'h4BFC] = 8'h00;
RAM[16'h4BFD] = 8'h00;
RAM[16'h4BFE] = 8'h00;
RAM[16'h4BFF] = 8'h00;
RAM[16'h4C00] = 8'h00;
RAM[16'h4C01] = 8'h00;
RAM[16'h4C02] = 8'h00;
RAM[16'h4C03] = 8'h00;
RAM[16'h4C04] = 8'h00;
RAM[16'h4C05] = 8'h00;
RAM[16'h4C06] = 8'h00;
RAM[16'h4C07] = 8'h00;
RAM[16'h4C08] = 8'h00;
RAM[16'h4C09] = 8'h00;
RAM[16'h4C0A] = 8'h00;
RAM[16'h4C0B] = 8'h00;
RAM[16'h4C0C] = 8'h00;
RAM[16'h4C0D] = 8'h00;
RAM[16'h4C0E] = 8'h00;
RAM[16'h4C0F] = 8'h00;
RAM[16'h4C10] = 8'h00;
RAM[16'h4C11] = 8'h00;
RAM[16'h4C12] = 8'h00;
RAM[16'h4C13] = 8'h00;
RAM[16'h4C14] = 8'h00;
RAM[16'h4C15] = 8'h00;
RAM[16'h4C16] = 8'h00;
RAM[16'h4C17] = 8'h00;
RAM[16'h4C18] = 8'h00;
RAM[16'h4C19] = 8'h00;
RAM[16'h4C1A] = 8'h00;
RAM[16'h4C1B] = 8'h00;
RAM[16'h4C1C] = 8'h00;
RAM[16'h4C1D] = 8'h00;
RAM[16'h4C1E] = 8'h00;
RAM[16'h4C1F] = 8'h00;
RAM[16'h4C20] = 8'h00;
RAM[16'h4C21] = 8'h00;
RAM[16'h4C22] = 8'h00;
RAM[16'h4C23] = 8'h00;
RAM[16'h4C24] = 8'h00;
RAM[16'h4C25] = 8'h00;
RAM[16'h4C26] = 8'h00;
RAM[16'h4C27] = 8'h00;
RAM[16'h4C28] = 8'h00;
RAM[16'h4C29] = 8'h00;
RAM[16'h4C2A] = 8'h00;
RAM[16'h4C2B] = 8'h00;
RAM[16'h4C2C] = 8'h00;
RAM[16'h4C2D] = 8'h00;
RAM[16'h4C2E] = 8'h00;
RAM[16'h4C2F] = 8'h00;
RAM[16'h4C30] = 8'h00;
RAM[16'h4C31] = 8'h00;
RAM[16'h4C32] = 8'h00;
RAM[16'h4C33] = 8'h00;
RAM[16'h4C34] = 8'h00;
RAM[16'h4C35] = 8'h00;
RAM[16'h4C36] = 8'h00;
RAM[16'h4C37] = 8'h00;
RAM[16'h4C38] = 8'h00;
RAM[16'h4C39] = 8'h00;
RAM[16'h4C3A] = 8'h00;
RAM[16'h4C3B] = 8'h00;
RAM[16'h4C3C] = 8'h00;
RAM[16'h4C3D] = 8'h00;
RAM[16'h4C3E] = 8'h00;
RAM[16'h4C3F] = 8'h00;
RAM[16'h4C40] = 8'h00;
RAM[16'h4C41] = 8'h00;
RAM[16'h4C42] = 8'h00;
RAM[16'h4C43] = 8'h00;
RAM[16'h4C44] = 8'h00;
RAM[16'h4C45] = 8'h00;
RAM[16'h4C46] = 8'h00;
RAM[16'h4C47] = 8'h00;
RAM[16'h4C48] = 8'h00;
RAM[16'h4C49] = 8'h00;
RAM[16'h4C4A] = 8'h00;
RAM[16'h4C4B] = 8'h00;
RAM[16'h4C4C] = 8'h00;
RAM[16'h4C4D] = 8'h00;
RAM[16'h4C4E] = 8'h00;
RAM[16'h4C4F] = 8'h00;
RAM[16'h4C50] = 8'h00;
RAM[16'h4C51] = 8'h00;
RAM[16'h4C52] = 8'h00;
RAM[16'h4C53] = 8'h00;
RAM[16'h4C54] = 8'h00;
RAM[16'h4C55] = 8'h00;
RAM[16'h4C56] = 8'h00;
RAM[16'h4C57] = 8'h00;
RAM[16'h4C58] = 8'h00;
RAM[16'h4C59] = 8'h00;
RAM[16'h4C5A] = 8'h00;
RAM[16'h4C5B] = 8'h00;
RAM[16'h4C5C] = 8'h00;
RAM[16'h4C5D] = 8'h00;
RAM[16'h4C5E] = 8'h00;
RAM[16'h4C5F] = 8'h00;
RAM[16'h4C60] = 8'h00;
RAM[16'h4C61] = 8'h00;
RAM[16'h4C62] = 8'h00;
RAM[16'h4C63] = 8'h00;
RAM[16'h4C64] = 8'h00;
RAM[16'h4C65] = 8'h00;
RAM[16'h4C66] = 8'h00;
RAM[16'h4C67] = 8'h00;
RAM[16'h4C68] = 8'h00;
RAM[16'h4C69] = 8'h00;
RAM[16'h4C6A] = 8'h00;
RAM[16'h4C6B] = 8'h00;
RAM[16'h4C6C] = 8'h00;
RAM[16'h4C6D] = 8'h00;
RAM[16'h4C6E] = 8'h00;
RAM[16'h4C6F] = 8'h00;
RAM[16'h4C70] = 8'h00;
RAM[16'h4C71] = 8'h00;
RAM[16'h4C72] = 8'h00;
RAM[16'h4C73] = 8'h00;
RAM[16'h4C74] = 8'h00;
RAM[16'h4C75] = 8'h00;
RAM[16'h4C76] = 8'h00;
RAM[16'h4C77] = 8'h00;
RAM[16'h4C78] = 8'h00;
RAM[16'h4C79] = 8'h00;
RAM[16'h4C7A] = 8'h00;
RAM[16'h4C7B] = 8'h00;
RAM[16'h4C7C] = 8'h00;
RAM[16'h4C7D] = 8'h00;
RAM[16'h4C7E] = 8'h00;
RAM[16'h4C7F] = 8'h00;
RAM[16'h4C80] = 8'h00;
RAM[16'h4C81] = 8'h00;
RAM[16'h4C82] = 8'h00;
RAM[16'h4C83] = 8'h00;
RAM[16'h4C84] = 8'h00;
RAM[16'h4C85] = 8'h00;
RAM[16'h4C86] = 8'h00;
RAM[16'h4C87] = 8'h00;
RAM[16'h4C88] = 8'h00;
RAM[16'h4C89] = 8'h00;
RAM[16'h4C8A] = 8'h00;
RAM[16'h4C8B] = 8'h00;
RAM[16'h4C8C] = 8'h00;
RAM[16'h4C8D] = 8'h00;
RAM[16'h4C8E] = 8'h00;
RAM[16'h4C8F] = 8'h00;
RAM[16'h4C90] = 8'h00;
RAM[16'h4C91] = 8'h00;
RAM[16'h4C92] = 8'h00;
RAM[16'h4C93] = 8'h00;
RAM[16'h4C94] = 8'h00;
RAM[16'h4C95] = 8'h00;
RAM[16'h4C96] = 8'h00;
RAM[16'h4C97] = 8'h00;
RAM[16'h4C98] = 8'h00;
RAM[16'h4C99] = 8'h00;
RAM[16'h4C9A] = 8'h00;
RAM[16'h4C9B] = 8'h00;
RAM[16'h4C9C] = 8'h00;
RAM[16'h4C9D] = 8'h00;
RAM[16'h4C9E] = 8'h00;
RAM[16'h4C9F] = 8'h00;
RAM[16'h4CA0] = 8'h00;
RAM[16'h4CA1] = 8'h00;
RAM[16'h4CA2] = 8'h00;
RAM[16'h4CA3] = 8'h00;
RAM[16'h4CA4] = 8'h00;
RAM[16'h4CA5] = 8'h00;
RAM[16'h4CA6] = 8'h00;
RAM[16'h4CA7] = 8'h00;
RAM[16'h4CA8] = 8'h00;
RAM[16'h4CA9] = 8'h00;
RAM[16'h4CAA] = 8'h00;
RAM[16'h4CAB] = 8'h00;
RAM[16'h4CAC] = 8'h00;
RAM[16'h4CAD] = 8'h00;
RAM[16'h4CAE] = 8'h00;
RAM[16'h4CAF] = 8'h00;
RAM[16'h4CB0] = 8'h00;
RAM[16'h4CB1] = 8'h00;
RAM[16'h4CB2] = 8'h00;
RAM[16'h4CB3] = 8'h00;
RAM[16'h4CB4] = 8'h00;
RAM[16'h4CB5] = 8'h00;
RAM[16'h4CB6] = 8'h00;
RAM[16'h4CB7] = 8'h00;
RAM[16'h4CB8] = 8'h00;
RAM[16'h4CB9] = 8'h00;
RAM[16'h4CBA] = 8'h00;
RAM[16'h4CBB] = 8'h00;
RAM[16'h4CBC] = 8'h00;
RAM[16'h4CBD] = 8'h00;
RAM[16'h4CBE] = 8'h00;
RAM[16'h4CBF] = 8'h00;
RAM[16'h4CC0] = 8'h00;
RAM[16'h4CC1] = 8'h00;
RAM[16'h4CC2] = 8'h00;
RAM[16'h4CC3] = 8'h00;
RAM[16'h4CC4] = 8'h00;
RAM[16'h4CC5] = 8'h00;
RAM[16'h4CC6] = 8'h00;
RAM[16'h4CC7] = 8'h00;
RAM[16'h4CC8] = 8'h00;
RAM[16'h4CC9] = 8'h00;
RAM[16'h4CCA] = 8'h00;
RAM[16'h4CCB] = 8'h00;
RAM[16'h4CCC] = 8'h00;
RAM[16'h4CCD] = 8'h00;
RAM[16'h4CCE] = 8'h00;
RAM[16'h4CCF] = 8'h00;
RAM[16'h4CD0] = 8'h00;
RAM[16'h4CD1] = 8'h00;
RAM[16'h4CD2] = 8'h00;
RAM[16'h4CD3] = 8'h00;
RAM[16'h4CD4] = 8'h00;
RAM[16'h4CD5] = 8'h00;
RAM[16'h4CD6] = 8'h00;
RAM[16'h4CD7] = 8'h00;
RAM[16'h4CD8] = 8'h00;
RAM[16'h4CD9] = 8'h00;
RAM[16'h4CDA] = 8'h00;
RAM[16'h4CDB] = 8'h00;
RAM[16'h4CDC] = 8'h00;
RAM[16'h4CDD] = 8'h00;
RAM[16'h4CDE] = 8'h00;
RAM[16'h4CDF] = 8'h00;
RAM[16'h4CE0] = 8'h00;
RAM[16'h4CE1] = 8'h00;
RAM[16'h4CE2] = 8'h00;
RAM[16'h4CE3] = 8'h00;
RAM[16'h4CE4] = 8'h00;
RAM[16'h4CE5] = 8'h00;
RAM[16'h4CE6] = 8'h00;
RAM[16'h4CE7] = 8'h00;
RAM[16'h4CE8] = 8'h00;
RAM[16'h4CE9] = 8'h00;
RAM[16'h4CEA] = 8'h00;
RAM[16'h4CEB] = 8'h00;
RAM[16'h4CEC] = 8'h00;
RAM[16'h4CED] = 8'h00;
RAM[16'h4CEE] = 8'h00;
RAM[16'h4CEF] = 8'h00;
RAM[16'h4CF0] = 8'h00;
RAM[16'h4CF1] = 8'h00;
RAM[16'h4CF2] = 8'h00;
RAM[16'h4CF3] = 8'h00;
RAM[16'h4CF4] = 8'h00;
RAM[16'h4CF5] = 8'h00;
RAM[16'h4CF6] = 8'h00;
RAM[16'h4CF7] = 8'h00;
RAM[16'h4CF8] = 8'h00;
RAM[16'h4CF9] = 8'h00;
RAM[16'h4CFA] = 8'h00;
RAM[16'h4CFB] = 8'h00;
RAM[16'h4CFC] = 8'h00;
RAM[16'h4CFD] = 8'h00;
RAM[16'h4CFE] = 8'h00;
RAM[16'h4CFF] = 8'h00;
RAM[16'h4D00] = 8'h00;
RAM[16'h4D01] = 8'h00;
RAM[16'h4D02] = 8'h00;
RAM[16'h4D03] = 8'h00;
RAM[16'h4D04] = 8'h00;
RAM[16'h4D05] = 8'h00;
RAM[16'h4D06] = 8'h00;
RAM[16'h4D07] = 8'h00;
RAM[16'h4D08] = 8'h00;
RAM[16'h4D09] = 8'h00;
RAM[16'h4D0A] = 8'h00;
RAM[16'h4D0B] = 8'h00;
RAM[16'h4D0C] = 8'h00;
RAM[16'h4D0D] = 8'h00;
RAM[16'h4D0E] = 8'h00;
RAM[16'h4D0F] = 8'h00;
RAM[16'h4D10] = 8'h00;
RAM[16'h4D11] = 8'h00;
RAM[16'h4D12] = 8'h00;
RAM[16'h4D13] = 8'h00;
RAM[16'h4D14] = 8'h00;
RAM[16'h4D15] = 8'h00;
RAM[16'h4D16] = 8'h00;
RAM[16'h4D17] = 8'h00;
RAM[16'h4D18] = 8'h00;
RAM[16'h4D19] = 8'h00;
RAM[16'h4D1A] = 8'h00;
RAM[16'h4D1B] = 8'h00;
RAM[16'h4D1C] = 8'h00;
RAM[16'h4D1D] = 8'h00;
RAM[16'h4D1E] = 8'h00;
RAM[16'h4D1F] = 8'h00;
RAM[16'h4D20] = 8'h00;
RAM[16'h4D21] = 8'h00;
RAM[16'h4D22] = 8'h00;
RAM[16'h4D23] = 8'h00;
RAM[16'h4D24] = 8'h00;
RAM[16'h4D25] = 8'h00;
RAM[16'h4D26] = 8'h00;
RAM[16'h4D27] = 8'h00;
RAM[16'h4D28] = 8'h00;
RAM[16'h4D29] = 8'h00;
RAM[16'h4D2A] = 8'h00;
RAM[16'h4D2B] = 8'h00;
RAM[16'h4D2C] = 8'h00;
RAM[16'h4D2D] = 8'h00;
RAM[16'h4D2E] = 8'h00;
RAM[16'h4D2F] = 8'h00;
RAM[16'h4D30] = 8'h00;
RAM[16'h4D31] = 8'h00;
RAM[16'h4D32] = 8'h00;
RAM[16'h4D33] = 8'h00;
RAM[16'h4D34] = 8'h00;
RAM[16'h4D35] = 8'h00;
RAM[16'h4D36] = 8'h00;
RAM[16'h4D37] = 8'h00;
RAM[16'h4D38] = 8'h00;
RAM[16'h4D39] = 8'h00;
RAM[16'h4D3A] = 8'h00;
RAM[16'h4D3B] = 8'h00;
RAM[16'h4D3C] = 8'h00;
RAM[16'h4D3D] = 8'h00;
RAM[16'h4D3E] = 8'h00;
RAM[16'h4D3F] = 8'h00;
RAM[16'h4D40] = 8'h00;
RAM[16'h4D41] = 8'h00;
RAM[16'h4D42] = 8'h00;
RAM[16'h4D43] = 8'h00;
RAM[16'h4D44] = 8'h00;
RAM[16'h4D45] = 8'h00;
RAM[16'h4D46] = 8'h00;
RAM[16'h4D47] = 8'h00;
RAM[16'h4D48] = 8'h00;
RAM[16'h4D49] = 8'h00;
RAM[16'h4D4A] = 8'h00;
RAM[16'h4D4B] = 8'h00;
RAM[16'h4D4C] = 8'h00;
RAM[16'h4D4D] = 8'h00;
RAM[16'h4D4E] = 8'h00;
RAM[16'h4D4F] = 8'h00;
RAM[16'h4D50] = 8'h00;
RAM[16'h4D51] = 8'h00;
RAM[16'h4D52] = 8'h00;
RAM[16'h4D53] = 8'h00;
RAM[16'h4D54] = 8'h00;
RAM[16'h4D55] = 8'h00;
RAM[16'h4D56] = 8'h00;
RAM[16'h4D57] = 8'h00;
RAM[16'h4D58] = 8'h00;
RAM[16'h4D59] = 8'h00;
RAM[16'h4D5A] = 8'h00;
RAM[16'h4D5B] = 8'h00;
RAM[16'h4D5C] = 8'h00;
RAM[16'h4D5D] = 8'h00;
RAM[16'h4D5E] = 8'h00;
RAM[16'h4D5F] = 8'h00;
RAM[16'h4D60] = 8'h00;
RAM[16'h4D61] = 8'h00;
RAM[16'h4D62] = 8'h00;
RAM[16'h4D63] = 8'h00;
RAM[16'h4D64] = 8'h00;
RAM[16'h4D65] = 8'h00;
RAM[16'h4D66] = 8'h00;
RAM[16'h4D67] = 8'h00;
RAM[16'h4D68] = 8'h00;
RAM[16'h4D69] = 8'h00;
RAM[16'h4D6A] = 8'h00;
RAM[16'h4D6B] = 8'h00;
RAM[16'h4D6C] = 8'h00;
RAM[16'h4D6D] = 8'h00;
RAM[16'h4D6E] = 8'h00;
RAM[16'h4D6F] = 8'h00;
RAM[16'h4D70] = 8'h00;
RAM[16'h4D71] = 8'h00;
RAM[16'h4D72] = 8'h00;
RAM[16'h4D73] = 8'h00;
RAM[16'h4D74] = 8'h00;
RAM[16'h4D75] = 8'h00;
RAM[16'h4D76] = 8'h00;
RAM[16'h4D77] = 8'h00;
RAM[16'h4D78] = 8'h00;
RAM[16'h4D79] = 8'h00;
RAM[16'h4D7A] = 8'h00;
RAM[16'h4D7B] = 8'h00;
RAM[16'h4D7C] = 8'h00;
RAM[16'h4D7D] = 8'h00;
RAM[16'h4D7E] = 8'h00;
RAM[16'h4D7F] = 8'h00;
RAM[16'h4D80] = 8'h00;
RAM[16'h4D81] = 8'h00;
RAM[16'h4D82] = 8'h00;
RAM[16'h4D83] = 8'h00;
RAM[16'h4D84] = 8'h00;
RAM[16'h4D85] = 8'h00;
RAM[16'h4D86] = 8'h00;
RAM[16'h4D87] = 8'h00;
RAM[16'h4D88] = 8'h00;
RAM[16'h4D89] = 8'h00;
RAM[16'h4D8A] = 8'h00;
RAM[16'h4D8B] = 8'h00;
RAM[16'h4D8C] = 8'h00;
RAM[16'h4D8D] = 8'h00;
RAM[16'h4D8E] = 8'h00;
RAM[16'h4D8F] = 8'h00;
RAM[16'h4D90] = 8'h00;
RAM[16'h4D91] = 8'h00;
RAM[16'h4D92] = 8'h00;
RAM[16'h4D93] = 8'h00;
RAM[16'h4D94] = 8'h00;
RAM[16'h4D95] = 8'h00;
RAM[16'h4D96] = 8'h00;
RAM[16'h4D97] = 8'h00;
RAM[16'h4D98] = 8'h00;
RAM[16'h4D99] = 8'h00;
RAM[16'h4D9A] = 8'h00;
RAM[16'h4D9B] = 8'h00;
RAM[16'h4D9C] = 8'h00;
RAM[16'h4D9D] = 8'h00;
RAM[16'h4D9E] = 8'h00;
RAM[16'h4D9F] = 8'h00;
RAM[16'h4DA0] = 8'h00;
RAM[16'h4DA1] = 8'h00;
RAM[16'h4DA2] = 8'h00;
RAM[16'h4DA3] = 8'h00;
RAM[16'h4DA4] = 8'h00;
RAM[16'h4DA5] = 8'h00;
RAM[16'h4DA6] = 8'h00;
RAM[16'h4DA7] = 8'h00;
RAM[16'h4DA8] = 8'h00;
RAM[16'h4DA9] = 8'h00;
RAM[16'h4DAA] = 8'h00;
RAM[16'h4DAB] = 8'h00;
RAM[16'h4DAC] = 8'h00;
RAM[16'h4DAD] = 8'h00;
RAM[16'h4DAE] = 8'h00;
RAM[16'h4DAF] = 8'h00;
RAM[16'h4DB0] = 8'h00;
RAM[16'h4DB1] = 8'h00;
RAM[16'h4DB2] = 8'h00;
RAM[16'h4DB3] = 8'h00;
RAM[16'h4DB4] = 8'h00;
RAM[16'h4DB5] = 8'h00;
RAM[16'h4DB6] = 8'h00;
RAM[16'h4DB7] = 8'h00;
RAM[16'h4DB8] = 8'h00;
RAM[16'h4DB9] = 8'h00;
RAM[16'h4DBA] = 8'h00;
RAM[16'h4DBB] = 8'h00;
RAM[16'h4DBC] = 8'h00;
RAM[16'h4DBD] = 8'h00;
RAM[16'h4DBE] = 8'h00;
RAM[16'h4DBF] = 8'h00;
RAM[16'h4DC0] = 8'h00;
RAM[16'h4DC1] = 8'h00;
RAM[16'h4DC2] = 8'h00;
RAM[16'h4DC3] = 8'h00;
RAM[16'h4DC4] = 8'h00;
RAM[16'h4DC5] = 8'h00;
RAM[16'h4DC6] = 8'h00;
RAM[16'h4DC7] = 8'h00;
RAM[16'h4DC8] = 8'h00;
RAM[16'h4DC9] = 8'h00;
RAM[16'h4DCA] = 8'h00;
RAM[16'h4DCB] = 8'h00;
RAM[16'h4DCC] = 8'h00;
RAM[16'h4DCD] = 8'h00;
RAM[16'h4DCE] = 8'h00;
RAM[16'h4DCF] = 8'h00;
RAM[16'h4DD0] = 8'h00;
RAM[16'h4DD1] = 8'h00;
RAM[16'h4DD2] = 8'h00;
RAM[16'h4DD3] = 8'h00;
RAM[16'h4DD4] = 8'h00;
RAM[16'h4DD5] = 8'h00;
RAM[16'h4DD6] = 8'h00;
RAM[16'h4DD7] = 8'h00;
RAM[16'h4DD8] = 8'h00;
RAM[16'h4DD9] = 8'h00;
RAM[16'h4DDA] = 8'h00;
RAM[16'h4DDB] = 8'h00;
RAM[16'h4DDC] = 8'h00;
RAM[16'h4DDD] = 8'h00;
RAM[16'h4DDE] = 8'h00;
RAM[16'h4DDF] = 8'h00;
RAM[16'h4DE0] = 8'h00;
RAM[16'h4DE1] = 8'h00;
RAM[16'h4DE2] = 8'h00;
RAM[16'h4DE3] = 8'h00;
RAM[16'h4DE4] = 8'h00;
RAM[16'h4DE5] = 8'h00;
RAM[16'h4DE6] = 8'h00;
RAM[16'h4DE7] = 8'h00;
RAM[16'h4DE8] = 8'h00;
RAM[16'h4DE9] = 8'h00;
RAM[16'h4DEA] = 8'h00;
RAM[16'h4DEB] = 8'h00;
RAM[16'h4DEC] = 8'h00;
RAM[16'h4DED] = 8'h00;
RAM[16'h4DEE] = 8'h00;
RAM[16'h4DEF] = 8'h00;
RAM[16'h4DF0] = 8'h00;
RAM[16'h4DF1] = 8'h00;
RAM[16'h4DF2] = 8'h00;
RAM[16'h4DF3] = 8'h00;
RAM[16'h4DF4] = 8'h00;
RAM[16'h4DF5] = 8'h00;
RAM[16'h4DF6] = 8'h00;
RAM[16'h4DF7] = 8'h00;
RAM[16'h4DF8] = 8'h00;
RAM[16'h4DF9] = 8'h00;
RAM[16'h4DFA] = 8'h00;
RAM[16'h4DFB] = 8'h00;
RAM[16'h4DFC] = 8'h00;
RAM[16'h4DFD] = 8'h00;
RAM[16'h4DFE] = 8'h00;
RAM[16'h4DFF] = 8'h00;
RAM[16'h4E00] = 8'h00;
RAM[16'h4E01] = 8'h00;
RAM[16'h4E02] = 8'h00;
RAM[16'h4E03] = 8'h00;
RAM[16'h4E04] = 8'h00;
RAM[16'h4E05] = 8'h00;
RAM[16'h4E06] = 8'h00;
RAM[16'h4E07] = 8'h00;
RAM[16'h4E08] = 8'h00;
RAM[16'h4E09] = 8'h00;
RAM[16'h4E0A] = 8'h00;
RAM[16'h4E0B] = 8'h00;
RAM[16'h4E0C] = 8'h00;
RAM[16'h4E0D] = 8'h00;
RAM[16'h4E0E] = 8'h00;
RAM[16'h4E0F] = 8'h00;
RAM[16'h4E10] = 8'h00;
RAM[16'h4E11] = 8'h00;
RAM[16'h4E12] = 8'h00;
RAM[16'h4E13] = 8'h00;
RAM[16'h4E14] = 8'h00;
RAM[16'h4E15] = 8'h00;
RAM[16'h4E16] = 8'h00;
RAM[16'h4E17] = 8'h00;
RAM[16'h4E18] = 8'h00;
RAM[16'h4E19] = 8'h00;
RAM[16'h4E1A] = 8'h00;
RAM[16'h4E1B] = 8'h00;
RAM[16'h4E1C] = 8'h00;
RAM[16'h4E1D] = 8'h00;
RAM[16'h4E1E] = 8'h00;
RAM[16'h4E1F] = 8'h00;
RAM[16'h4E20] = 8'h00;
RAM[16'h4E21] = 8'h00;
RAM[16'h4E22] = 8'h00;
RAM[16'h4E23] = 8'h00;
RAM[16'h4E24] = 8'h00;
RAM[16'h4E25] = 8'h00;
RAM[16'h4E26] = 8'h00;
RAM[16'h4E27] = 8'h00;
RAM[16'h4E28] = 8'h00;
RAM[16'h4E29] = 8'h00;
RAM[16'h4E2A] = 8'h00;
RAM[16'h4E2B] = 8'h00;
RAM[16'h4E2C] = 8'h00;
RAM[16'h4E2D] = 8'h00;
RAM[16'h4E2E] = 8'h00;
RAM[16'h4E2F] = 8'h00;
RAM[16'h4E30] = 8'h00;
RAM[16'h4E31] = 8'h00;
RAM[16'h4E32] = 8'h00;
RAM[16'h4E33] = 8'h00;
RAM[16'h4E34] = 8'h00;
RAM[16'h4E35] = 8'h00;
RAM[16'h4E36] = 8'h00;
RAM[16'h4E37] = 8'h00;
RAM[16'h4E38] = 8'h00;
RAM[16'h4E39] = 8'h00;
RAM[16'h4E3A] = 8'h00;
RAM[16'h4E3B] = 8'h00;
RAM[16'h4E3C] = 8'h00;
RAM[16'h4E3D] = 8'h00;
RAM[16'h4E3E] = 8'h00;
RAM[16'h4E3F] = 8'h00;
RAM[16'h4E40] = 8'h00;
RAM[16'h4E41] = 8'h00;
RAM[16'h4E42] = 8'h00;
RAM[16'h4E43] = 8'h00;
RAM[16'h4E44] = 8'h00;
RAM[16'h4E45] = 8'h00;
RAM[16'h4E46] = 8'h00;
RAM[16'h4E47] = 8'h00;
RAM[16'h4E48] = 8'h00;
RAM[16'h4E49] = 8'h00;
RAM[16'h4E4A] = 8'h00;
RAM[16'h4E4B] = 8'h00;
RAM[16'h4E4C] = 8'h00;
RAM[16'h4E4D] = 8'h00;
RAM[16'h4E4E] = 8'h00;
RAM[16'h4E4F] = 8'h00;
RAM[16'h4E50] = 8'h00;
RAM[16'h4E51] = 8'h00;
RAM[16'h4E52] = 8'h00;
RAM[16'h4E53] = 8'h00;
RAM[16'h4E54] = 8'h00;
RAM[16'h4E55] = 8'h00;
RAM[16'h4E56] = 8'h00;
RAM[16'h4E57] = 8'h00;
RAM[16'h4E58] = 8'h00;
RAM[16'h4E59] = 8'h00;
RAM[16'h4E5A] = 8'h00;
RAM[16'h4E5B] = 8'h00;
RAM[16'h4E5C] = 8'h00;
RAM[16'h4E5D] = 8'h00;
RAM[16'h4E5E] = 8'h00;
RAM[16'h4E5F] = 8'h00;
RAM[16'h4E60] = 8'h00;
RAM[16'h4E61] = 8'h00;
RAM[16'h4E62] = 8'h00;
RAM[16'h4E63] = 8'h00;
RAM[16'h4E64] = 8'h00;
RAM[16'h4E65] = 8'h00;
RAM[16'h4E66] = 8'h00;
RAM[16'h4E67] = 8'h00;
RAM[16'h4E68] = 8'h00;
RAM[16'h4E69] = 8'h00;
RAM[16'h4E6A] = 8'h00;
RAM[16'h4E6B] = 8'h00;
RAM[16'h4E6C] = 8'h00;
RAM[16'h4E6D] = 8'h00;
RAM[16'h4E6E] = 8'h00;
RAM[16'h4E6F] = 8'h00;
RAM[16'h4E70] = 8'h00;
RAM[16'h4E71] = 8'h00;
RAM[16'h4E72] = 8'h00;
RAM[16'h4E73] = 8'h00;
RAM[16'h4E74] = 8'h00;
RAM[16'h4E75] = 8'h00;
RAM[16'h4E76] = 8'h00;
RAM[16'h4E77] = 8'h00;
RAM[16'h4E78] = 8'h00;
RAM[16'h4E79] = 8'h00;
RAM[16'h4E7A] = 8'h00;
RAM[16'h4E7B] = 8'h00;
RAM[16'h4E7C] = 8'h00;
RAM[16'h4E7D] = 8'h00;
RAM[16'h4E7E] = 8'h00;
RAM[16'h4E7F] = 8'h00;
RAM[16'h4E80] = 8'h00;
RAM[16'h4E81] = 8'h00;
RAM[16'h4E82] = 8'h00;
RAM[16'h4E83] = 8'h00;
RAM[16'h4E84] = 8'h00;
RAM[16'h4E85] = 8'h00;
RAM[16'h4E86] = 8'h00;
RAM[16'h4E87] = 8'h00;
RAM[16'h4E88] = 8'h00;
RAM[16'h4E89] = 8'h00;
RAM[16'h4E8A] = 8'h00;
RAM[16'h4E8B] = 8'h00;
RAM[16'h4E8C] = 8'h00;
RAM[16'h4E8D] = 8'h00;
RAM[16'h4E8E] = 8'h00;
RAM[16'h4E8F] = 8'h00;
RAM[16'h4E90] = 8'h00;
RAM[16'h4E91] = 8'h00;
RAM[16'h4E92] = 8'h00;
RAM[16'h4E93] = 8'h00;
RAM[16'h4E94] = 8'h00;
RAM[16'h4E95] = 8'h00;
RAM[16'h4E96] = 8'h00;
RAM[16'h4E97] = 8'h00;
RAM[16'h4E98] = 8'h00;
RAM[16'h4E99] = 8'h00;
RAM[16'h4E9A] = 8'h00;
RAM[16'h4E9B] = 8'h00;
RAM[16'h4E9C] = 8'h00;
RAM[16'h4E9D] = 8'h00;
RAM[16'h4E9E] = 8'h00;
RAM[16'h4E9F] = 8'h00;
RAM[16'h4EA0] = 8'h00;
RAM[16'h4EA1] = 8'h00;
RAM[16'h4EA2] = 8'h00;
RAM[16'h4EA3] = 8'h00;
RAM[16'h4EA4] = 8'h00;
RAM[16'h4EA5] = 8'h00;
RAM[16'h4EA6] = 8'h00;
RAM[16'h4EA7] = 8'h00;
RAM[16'h4EA8] = 8'h00;
RAM[16'h4EA9] = 8'h00;
RAM[16'h4EAA] = 8'h00;
RAM[16'h4EAB] = 8'h00;
RAM[16'h4EAC] = 8'h00;
RAM[16'h4EAD] = 8'h00;
RAM[16'h4EAE] = 8'h00;
RAM[16'h4EAF] = 8'h00;
RAM[16'h4EB0] = 8'h00;
RAM[16'h4EB1] = 8'h00;
RAM[16'h4EB2] = 8'h00;
RAM[16'h4EB3] = 8'h00;
RAM[16'h4EB4] = 8'h00;
RAM[16'h4EB5] = 8'h00;
RAM[16'h4EB6] = 8'h00;
RAM[16'h4EB7] = 8'h00;
RAM[16'h4EB8] = 8'h00;
RAM[16'h4EB9] = 8'h00;
RAM[16'h4EBA] = 8'h00;
RAM[16'h4EBB] = 8'h00;
RAM[16'h4EBC] = 8'h00;
RAM[16'h4EBD] = 8'h00;
RAM[16'h4EBE] = 8'h00;
RAM[16'h4EBF] = 8'h00;
RAM[16'h4EC0] = 8'h00;
RAM[16'h4EC1] = 8'h00;
RAM[16'h4EC2] = 8'h00;
RAM[16'h4EC3] = 8'h00;
RAM[16'h4EC4] = 8'h00;
RAM[16'h4EC5] = 8'h00;
RAM[16'h4EC6] = 8'h00;
RAM[16'h4EC7] = 8'h00;
RAM[16'h4EC8] = 8'h00;
RAM[16'h4EC9] = 8'h00;
RAM[16'h4ECA] = 8'h00;
RAM[16'h4ECB] = 8'h00;
RAM[16'h4ECC] = 8'h00;
RAM[16'h4ECD] = 8'h00;
RAM[16'h4ECE] = 8'h00;
RAM[16'h4ECF] = 8'h00;
RAM[16'h4ED0] = 8'h00;
RAM[16'h4ED1] = 8'h00;
RAM[16'h4ED2] = 8'h00;
RAM[16'h4ED3] = 8'h00;
RAM[16'h4ED4] = 8'h00;
RAM[16'h4ED5] = 8'h00;
RAM[16'h4ED6] = 8'h00;
RAM[16'h4ED7] = 8'h00;
RAM[16'h4ED8] = 8'h00;
RAM[16'h4ED9] = 8'h00;
RAM[16'h4EDA] = 8'h00;
RAM[16'h4EDB] = 8'h00;
RAM[16'h4EDC] = 8'h00;
RAM[16'h4EDD] = 8'h00;
RAM[16'h4EDE] = 8'h00;
RAM[16'h4EDF] = 8'h00;
RAM[16'h4EE0] = 8'h00;
RAM[16'h4EE1] = 8'h00;
RAM[16'h4EE2] = 8'h00;
RAM[16'h4EE3] = 8'h00;
RAM[16'h4EE4] = 8'h00;
RAM[16'h4EE5] = 8'h00;
RAM[16'h4EE6] = 8'h00;
RAM[16'h4EE7] = 8'h00;
RAM[16'h4EE8] = 8'h00;
RAM[16'h4EE9] = 8'h00;
RAM[16'h4EEA] = 8'h00;
RAM[16'h4EEB] = 8'h00;
RAM[16'h4EEC] = 8'h00;
RAM[16'h4EED] = 8'h00;
RAM[16'h4EEE] = 8'h00;
RAM[16'h4EEF] = 8'h00;
RAM[16'h4EF0] = 8'h00;
RAM[16'h4EF1] = 8'h00;
RAM[16'h4EF2] = 8'h00;
RAM[16'h4EF3] = 8'h00;
RAM[16'h4EF4] = 8'h00;
RAM[16'h4EF5] = 8'h00;
RAM[16'h4EF6] = 8'h00;
RAM[16'h4EF7] = 8'h00;
RAM[16'h4EF8] = 8'h00;
RAM[16'h4EF9] = 8'h00;
RAM[16'h4EFA] = 8'h00;
RAM[16'h4EFB] = 8'h00;
RAM[16'h4EFC] = 8'h00;
RAM[16'h4EFD] = 8'h00;
RAM[16'h4EFE] = 8'h00;
RAM[16'h4EFF] = 8'h00;
RAM[16'h4F00] = 8'h00;
RAM[16'h4F01] = 8'h00;
RAM[16'h4F02] = 8'h00;
RAM[16'h4F03] = 8'h00;
RAM[16'h4F04] = 8'h00;
RAM[16'h4F05] = 8'h00;
RAM[16'h4F06] = 8'h00;
RAM[16'h4F07] = 8'h00;
RAM[16'h4F08] = 8'h00;
RAM[16'h4F09] = 8'h00;
RAM[16'h4F0A] = 8'h00;
RAM[16'h4F0B] = 8'h00;
RAM[16'h4F0C] = 8'h00;
RAM[16'h4F0D] = 8'h00;
RAM[16'h4F0E] = 8'h00;
RAM[16'h4F0F] = 8'h00;
RAM[16'h4F10] = 8'h00;
RAM[16'h4F11] = 8'h00;
RAM[16'h4F12] = 8'h00;
RAM[16'h4F13] = 8'h00;
RAM[16'h4F14] = 8'h00;
RAM[16'h4F15] = 8'h00;
RAM[16'h4F16] = 8'h00;
RAM[16'h4F17] = 8'h00;
RAM[16'h4F18] = 8'h00;
RAM[16'h4F19] = 8'h00;
RAM[16'h4F1A] = 8'h00;
RAM[16'h4F1B] = 8'h00;
RAM[16'h4F1C] = 8'h00;
RAM[16'h4F1D] = 8'h00;
RAM[16'h4F1E] = 8'h00;
RAM[16'h4F1F] = 8'h00;
RAM[16'h4F20] = 8'h00;
RAM[16'h4F21] = 8'h00;
RAM[16'h4F22] = 8'h00;
RAM[16'h4F23] = 8'h00;
RAM[16'h4F24] = 8'h00;
RAM[16'h4F25] = 8'h00;
RAM[16'h4F26] = 8'h00;
RAM[16'h4F27] = 8'h00;
RAM[16'h4F28] = 8'h00;
RAM[16'h4F29] = 8'h00;
RAM[16'h4F2A] = 8'h00;
RAM[16'h4F2B] = 8'h00;
RAM[16'h4F2C] = 8'h00;
RAM[16'h4F2D] = 8'h00;
RAM[16'h4F2E] = 8'h00;
RAM[16'h4F2F] = 8'h00;
RAM[16'h4F30] = 8'h00;
RAM[16'h4F31] = 8'h00;
RAM[16'h4F32] = 8'h00;
RAM[16'h4F33] = 8'h00;
RAM[16'h4F34] = 8'h00;
RAM[16'h4F35] = 8'h00;
RAM[16'h4F36] = 8'h00;
RAM[16'h4F37] = 8'h00;
RAM[16'h4F38] = 8'h00;
RAM[16'h4F39] = 8'h00;
RAM[16'h4F3A] = 8'h00;
RAM[16'h4F3B] = 8'h00;
RAM[16'h4F3C] = 8'h00;
RAM[16'h4F3D] = 8'h00;
RAM[16'h4F3E] = 8'h00;
RAM[16'h4F3F] = 8'h00;
RAM[16'h4F40] = 8'h00;
RAM[16'h4F41] = 8'h00;
RAM[16'h4F42] = 8'h00;
RAM[16'h4F43] = 8'h00;
RAM[16'h4F44] = 8'h00;
RAM[16'h4F45] = 8'h00;
RAM[16'h4F46] = 8'h00;
RAM[16'h4F47] = 8'h00;
RAM[16'h4F48] = 8'h00;
RAM[16'h4F49] = 8'h00;
RAM[16'h4F4A] = 8'h00;
RAM[16'h4F4B] = 8'h00;
RAM[16'h4F4C] = 8'h00;
RAM[16'h4F4D] = 8'h00;
RAM[16'h4F4E] = 8'h00;
RAM[16'h4F4F] = 8'h00;
RAM[16'h4F50] = 8'h00;
RAM[16'h4F51] = 8'h00;
RAM[16'h4F52] = 8'h00;
RAM[16'h4F53] = 8'h00;
RAM[16'h4F54] = 8'h00;
RAM[16'h4F55] = 8'h00;
RAM[16'h4F56] = 8'h00;
RAM[16'h4F57] = 8'h00;
RAM[16'h4F58] = 8'h00;
RAM[16'h4F59] = 8'h00;
RAM[16'h4F5A] = 8'h00;
RAM[16'h4F5B] = 8'h00;
RAM[16'h4F5C] = 8'h00;
RAM[16'h4F5D] = 8'h00;
RAM[16'h4F5E] = 8'h00;
RAM[16'h4F5F] = 8'h00;
RAM[16'h4F60] = 8'h00;
RAM[16'h4F61] = 8'h00;
RAM[16'h4F62] = 8'h00;
RAM[16'h4F63] = 8'h00;
RAM[16'h4F64] = 8'h00;
RAM[16'h4F65] = 8'h00;
RAM[16'h4F66] = 8'h00;
RAM[16'h4F67] = 8'h00;
RAM[16'h4F68] = 8'h00;
RAM[16'h4F69] = 8'h00;
RAM[16'h4F6A] = 8'h00;
RAM[16'h4F6B] = 8'h00;
RAM[16'h4F6C] = 8'h00;
RAM[16'h4F6D] = 8'h00;
RAM[16'h4F6E] = 8'h00;
RAM[16'h4F6F] = 8'h00;
RAM[16'h4F70] = 8'h00;
RAM[16'h4F71] = 8'h00;
RAM[16'h4F72] = 8'h00;
RAM[16'h4F73] = 8'h00;
RAM[16'h4F74] = 8'h00;
RAM[16'h4F75] = 8'h00;
RAM[16'h4F76] = 8'h00;
RAM[16'h4F77] = 8'h00;
RAM[16'h4F78] = 8'h00;
RAM[16'h4F79] = 8'h00;
RAM[16'h4F7A] = 8'h00;
RAM[16'h4F7B] = 8'h00;
RAM[16'h4F7C] = 8'h00;
RAM[16'h4F7D] = 8'h00;
RAM[16'h4F7E] = 8'h00;
RAM[16'h4F7F] = 8'h00;
RAM[16'h4F80] = 8'h00;
RAM[16'h4F81] = 8'h00;
RAM[16'h4F82] = 8'h00;
RAM[16'h4F83] = 8'h00;
RAM[16'h4F84] = 8'h00;
RAM[16'h4F85] = 8'h00;
RAM[16'h4F86] = 8'h00;
RAM[16'h4F87] = 8'h00;
RAM[16'h4F88] = 8'h00;
RAM[16'h4F89] = 8'h00;
RAM[16'h4F8A] = 8'h00;
RAM[16'h4F8B] = 8'h00;
RAM[16'h4F8C] = 8'h00;
RAM[16'h4F8D] = 8'h00;
RAM[16'h4F8E] = 8'h00;
RAM[16'h4F8F] = 8'h00;
RAM[16'h4F90] = 8'h00;
RAM[16'h4F91] = 8'h00;
RAM[16'h4F92] = 8'h00;
RAM[16'h4F93] = 8'h00;
RAM[16'h4F94] = 8'h00;
RAM[16'h4F95] = 8'h00;
RAM[16'h4F96] = 8'h00;
RAM[16'h4F97] = 8'h00;
RAM[16'h4F98] = 8'h00;
RAM[16'h4F99] = 8'h00;
RAM[16'h4F9A] = 8'h00;
RAM[16'h4F9B] = 8'h00;
RAM[16'h4F9C] = 8'h00;
RAM[16'h4F9D] = 8'h00;
RAM[16'h4F9E] = 8'h00;
RAM[16'h4F9F] = 8'h00;
RAM[16'h4FA0] = 8'h00;
RAM[16'h4FA1] = 8'h00;
RAM[16'h4FA2] = 8'h00;
RAM[16'h4FA3] = 8'h00;
RAM[16'h4FA4] = 8'h00;
RAM[16'h4FA5] = 8'h00;
RAM[16'h4FA6] = 8'h00;
RAM[16'h4FA7] = 8'h00;
RAM[16'h4FA8] = 8'h00;
RAM[16'h4FA9] = 8'h00;
RAM[16'h4FAA] = 8'h00;
RAM[16'h4FAB] = 8'h00;
RAM[16'h4FAC] = 8'h00;
RAM[16'h4FAD] = 8'h00;
RAM[16'h4FAE] = 8'h00;
RAM[16'h4FAF] = 8'h00;
RAM[16'h4FB0] = 8'h00;
RAM[16'h4FB1] = 8'h00;
RAM[16'h4FB2] = 8'h00;
RAM[16'h4FB3] = 8'h00;
RAM[16'h4FB4] = 8'h00;
RAM[16'h4FB5] = 8'h00;
RAM[16'h4FB6] = 8'h00;
RAM[16'h4FB7] = 8'h00;
RAM[16'h4FB8] = 8'h00;
RAM[16'h4FB9] = 8'h00;
RAM[16'h4FBA] = 8'h00;
RAM[16'h4FBB] = 8'h00;
RAM[16'h4FBC] = 8'h00;
RAM[16'h4FBD] = 8'h00;
RAM[16'h4FBE] = 8'h00;
RAM[16'h4FBF] = 8'h00;
RAM[16'h4FC0] = 8'h00;
RAM[16'h4FC1] = 8'h00;
RAM[16'h4FC2] = 8'h00;
RAM[16'h4FC3] = 8'h00;
RAM[16'h4FC4] = 8'h00;
RAM[16'h4FC5] = 8'h00;
RAM[16'h4FC6] = 8'h00;
RAM[16'h4FC7] = 8'h00;
RAM[16'h4FC8] = 8'h00;
RAM[16'h4FC9] = 8'h00;
RAM[16'h4FCA] = 8'h00;
RAM[16'h4FCB] = 8'h00;
RAM[16'h4FCC] = 8'h00;
RAM[16'h4FCD] = 8'h00;
RAM[16'h4FCE] = 8'h00;
RAM[16'h4FCF] = 8'h00;
RAM[16'h4FD0] = 8'h00;
RAM[16'h4FD1] = 8'h00;
RAM[16'h4FD2] = 8'h00;
RAM[16'h4FD3] = 8'h00;
RAM[16'h4FD4] = 8'h00;
RAM[16'h4FD5] = 8'h00;
RAM[16'h4FD6] = 8'h00;
RAM[16'h4FD7] = 8'h00;
RAM[16'h4FD8] = 8'h00;
RAM[16'h4FD9] = 8'h00;
RAM[16'h4FDA] = 8'h00;
RAM[16'h4FDB] = 8'h00;
RAM[16'h4FDC] = 8'h00;
RAM[16'h4FDD] = 8'h00;
RAM[16'h4FDE] = 8'h00;
RAM[16'h4FDF] = 8'h00;
RAM[16'h4FE0] = 8'h00;
RAM[16'h4FE1] = 8'h00;
RAM[16'h4FE2] = 8'h00;
RAM[16'h4FE3] = 8'h00;
RAM[16'h4FE4] = 8'h00;
RAM[16'h4FE5] = 8'h00;
RAM[16'h4FE6] = 8'h00;
RAM[16'h4FE7] = 8'h00;
RAM[16'h4FE8] = 8'h00;
RAM[16'h4FE9] = 8'h00;
RAM[16'h4FEA] = 8'h00;
RAM[16'h4FEB] = 8'h00;
RAM[16'h4FEC] = 8'h00;
RAM[16'h4FED] = 8'h00;
RAM[16'h4FEE] = 8'h00;
RAM[16'h4FEF] = 8'h00;
RAM[16'h4FF0] = 8'h00;
RAM[16'h4FF1] = 8'h00;
RAM[16'h4FF2] = 8'h00;
RAM[16'h4FF3] = 8'h00;
RAM[16'h4FF4] = 8'h00;
RAM[16'h4FF5] = 8'h00;
RAM[16'h4FF6] = 8'h00;
RAM[16'h4FF7] = 8'h00;
RAM[16'h4FF8] = 8'h00;
RAM[16'h4FF9] = 8'h00;
RAM[16'h4FFA] = 8'h00;
RAM[16'h4FFB] = 8'h00;
RAM[16'h4FFC] = 8'h00;
RAM[16'h4FFD] = 8'h00;
RAM[16'h4FFE] = 8'h00;
RAM[16'h4FFF] = 8'h00;
RAM[16'h5000] = 8'h00;
RAM[16'h5001] = 8'h00;
RAM[16'h5002] = 8'h00;
RAM[16'h5003] = 8'h00;
RAM[16'h5004] = 8'h00;
RAM[16'h5005] = 8'h00;
RAM[16'h5006] = 8'h00;
RAM[16'h5007] = 8'h00;
RAM[16'h5008] = 8'h00;
RAM[16'h5009] = 8'h00;
RAM[16'h500A] = 8'h00;
RAM[16'h500B] = 8'h00;
RAM[16'h500C] = 8'h00;
RAM[16'h500D] = 8'h00;
RAM[16'h500E] = 8'h00;
RAM[16'h500F] = 8'h00;
RAM[16'h5010] = 8'h00;
RAM[16'h5011] = 8'h00;
RAM[16'h5012] = 8'h00;
RAM[16'h5013] = 8'h00;
RAM[16'h5014] = 8'h00;
RAM[16'h5015] = 8'h00;
RAM[16'h5016] = 8'h00;
RAM[16'h5017] = 8'h00;
RAM[16'h5018] = 8'h00;
RAM[16'h5019] = 8'h00;
RAM[16'h501A] = 8'h00;
RAM[16'h501B] = 8'h00;
RAM[16'h501C] = 8'h00;
RAM[16'h501D] = 8'h00;
RAM[16'h501E] = 8'h00;
RAM[16'h501F] = 8'h00;
RAM[16'h5020] = 8'h00;
RAM[16'h5021] = 8'h00;
RAM[16'h5022] = 8'h00;
RAM[16'h5023] = 8'h00;
RAM[16'h5024] = 8'h00;
RAM[16'h5025] = 8'h00;
RAM[16'h5026] = 8'h00;
RAM[16'h5027] = 8'h00;
RAM[16'h5028] = 8'h00;
RAM[16'h5029] = 8'h00;
RAM[16'h502A] = 8'h00;
RAM[16'h502B] = 8'h00;
RAM[16'h502C] = 8'h00;
RAM[16'h502D] = 8'h00;
RAM[16'h502E] = 8'h00;
RAM[16'h502F] = 8'h00;
RAM[16'h5030] = 8'h00;
RAM[16'h5031] = 8'h00;
RAM[16'h5032] = 8'h00;
RAM[16'h5033] = 8'h00;
RAM[16'h5034] = 8'h00;
RAM[16'h5035] = 8'h00;
RAM[16'h5036] = 8'h00;
RAM[16'h5037] = 8'h00;
RAM[16'h5038] = 8'h00;
RAM[16'h5039] = 8'h00;
RAM[16'h503A] = 8'h00;
RAM[16'h503B] = 8'h00;
RAM[16'h503C] = 8'h00;
RAM[16'h503D] = 8'h00;
RAM[16'h503E] = 8'h00;
RAM[16'h503F] = 8'h00;
RAM[16'h5040] = 8'h00;
RAM[16'h5041] = 8'h00;
RAM[16'h5042] = 8'h00;
RAM[16'h5043] = 8'h00;
RAM[16'h5044] = 8'h00;
RAM[16'h5045] = 8'h00;
RAM[16'h5046] = 8'h00;
RAM[16'h5047] = 8'h00;
RAM[16'h5048] = 8'h00;
RAM[16'h5049] = 8'h00;
RAM[16'h504A] = 8'h00;
RAM[16'h504B] = 8'h00;
RAM[16'h504C] = 8'h00;
RAM[16'h504D] = 8'h00;
RAM[16'h504E] = 8'h00;
RAM[16'h504F] = 8'h00;
RAM[16'h5050] = 8'h00;
RAM[16'h5051] = 8'h00;
RAM[16'h5052] = 8'h00;
RAM[16'h5053] = 8'h00;
RAM[16'h5054] = 8'h00;
RAM[16'h5055] = 8'h00;
RAM[16'h5056] = 8'h00;
RAM[16'h5057] = 8'h00;
RAM[16'h5058] = 8'h00;
RAM[16'h5059] = 8'h00;
RAM[16'h505A] = 8'h00;
RAM[16'h505B] = 8'h00;
RAM[16'h505C] = 8'h00;
RAM[16'h505D] = 8'h00;
RAM[16'h505E] = 8'h00;
RAM[16'h505F] = 8'h00;
RAM[16'h5060] = 8'h00;
RAM[16'h5061] = 8'h00;
RAM[16'h5062] = 8'h00;
RAM[16'h5063] = 8'h00;
RAM[16'h5064] = 8'h00;
RAM[16'h5065] = 8'h00;
RAM[16'h5066] = 8'h00;
RAM[16'h5067] = 8'h00;
RAM[16'h5068] = 8'h00;
RAM[16'h5069] = 8'h00;
RAM[16'h506A] = 8'h00;
RAM[16'h506B] = 8'h00;
RAM[16'h506C] = 8'h00;
RAM[16'h506D] = 8'h00;
RAM[16'h506E] = 8'h00;
RAM[16'h506F] = 8'h00;
RAM[16'h5070] = 8'h00;
RAM[16'h5071] = 8'h00;
RAM[16'h5072] = 8'h00;
RAM[16'h5073] = 8'h00;
RAM[16'h5074] = 8'h00;
RAM[16'h5075] = 8'h00;
RAM[16'h5076] = 8'h00;
RAM[16'h5077] = 8'h00;
RAM[16'h5078] = 8'h00;
RAM[16'h5079] = 8'h00;
RAM[16'h507A] = 8'h00;
RAM[16'h507B] = 8'h00;
RAM[16'h507C] = 8'h00;
RAM[16'h507D] = 8'h00;
RAM[16'h507E] = 8'h00;
RAM[16'h507F] = 8'h00;
RAM[16'h5080] = 8'h00;
RAM[16'h5081] = 8'h00;
RAM[16'h5082] = 8'h00;
RAM[16'h5083] = 8'h00;
RAM[16'h5084] = 8'h00;
RAM[16'h5085] = 8'h00;
RAM[16'h5086] = 8'h00;
RAM[16'h5087] = 8'h00;
RAM[16'h5088] = 8'h00;
RAM[16'h5089] = 8'h00;
RAM[16'h508A] = 8'h00;
RAM[16'h508B] = 8'h00;
RAM[16'h508C] = 8'h00;
RAM[16'h508D] = 8'h00;
RAM[16'h508E] = 8'h00;
RAM[16'h508F] = 8'h00;
RAM[16'h5090] = 8'h00;
RAM[16'h5091] = 8'h00;
RAM[16'h5092] = 8'h00;
RAM[16'h5093] = 8'h00;
RAM[16'h5094] = 8'h00;
RAM[16'h5095] = 8'h00;
RAM[16'h5096] = 8'h00;
RAM[16'h5097] = 8'h00;
RAM[16'h5098] = 8'h00;
RAM[16'h5099] = 8'h00;
RAM[16'h509A] = 8'h00;
RAM[16'h509B] = 8'h00;
RAM[16'h509C] = 8'h00;
RAM[16'h509D] = 8'h00;
RAM[16'h509E] = 8'h00;
RAM[16'h509F] = 8'h00;
RAM[16'h50A0] = 8'h00;
RAM[16'h50A1] = 8'h00;
RAM[16'h50A2] = 8'h00;
RAM[16'h50A3] = 8'h00;
RAM[16'h50A4] = 8'h00;
RAM[16'h50A5] = 8'h00;
RAM[16'h50A6] = 8'h00;
RAM[16'h50A7] = 8'h00;
RAM[16'h50A8] = 8'h00;
RAM[16'h50A9] = 8'h00;
RAM[16'h50AA] = 8'h00;
RAM[16'h50AB] = 8'h00;
RAM[16'h50AC] = 8'h00;
RAM[16'h50AD] = 8'h00;
RAM[16'h50AE] = 8'h00;
RAM[16'h50AF] = 8'h00;
RAM[16'h50B0] = 8'h00;
RAM[16'h50B1] = 8'h00;
RAM[16'h50B2] = 8'h00;
RAM[16'h50B3] = 8'h00;
RAM[16'h50B4] = 8'h00;
RAM[16'h50B5] = 8'h00;
RAM[16'h50B6] = 8'h00;
RAM[16'h50B7] = 8'h00;
RAM[16'h50B8] = 8'h00;
RAM[16'h50B9] = 8'h00;
RAM[16'h50BA] = 8'h00;
RAM[16'h50BB] = 8'h00;
RAM[16'h50BC] = 8'h00;
RAM[16'h50BD] = 8'h00;
RAM[16'h50BE] = 8'h00;
RAM[16'h50BF] = 8'h00;
RAM[16'h50C0] = 8'h00;
RAM[16'h50C1] = 8'h00;
RAM[16'h50C2] = 8'h00;
RAM[16'h50C3] = 8'h00;
RAM[16'h50C4] = 8'h00;
RAM[16'h50C5] = 8'h00;
RAM[16'h50C6] = 8'h00;
RAM[16'h50C7] = 8'h00;
RAM[16'h50C8] = 8'h00;
RAM[16'h50C9] = 8'h00;
RAM[16'h50CA] = 8'h00;
RAM[16'h50CB] = 8'h00;
RAM[16'h50CC] = 8'h00;
RAM[16'h50CD] = 8'h00;
RAM[16'h50CE] = 8'h00;
RAM[16'h50CF] = 8'h00;
RAM[16'h50D0] = 8'h00;
RAM[16'h50D1] = 8'h00;
RAM[16'h50D2] = 8'h00;
RAM[16'h50D3] = 8'h00;
RAM[16'h50D4] = 8'h00;
RAM[16'h50D5] = 8'h00;
RAM[16'h50D6] = 8'h00;
RAM[16'h50D7] = 8'h00;
RAM[16'h50D8] = 8'h00;
RAM[16'h50D9] = 8'h00;
RAM[16'h50DA] = 8'h00;
RAM[16'h50DB] = 8'h00;
RAM[16'h50DC] = 8'h00;
RAM[16'h50DD] = 8'h00;
RAM[16'h50DE] = 8'h00;
RAM[16'h50DF] = 8'h00;
RAM[16'h50E0] = 8'h00;
RAM[16'h50E1] = 8'h00;
RAM[16'h50E2] = 8'h00;
RAM[16'h50E3] = 8'h00;
RAM[16'h50E4] = 8'h00;
RAM[16'h50E5] = 8'h00;
RAM[16'h50E6] = 8'h00;
RAM[16'h50E7] = 8'h00;
RAM[16'h50E8] = 8'h00;
RAM[16'h50E9] = 8'h00;
RAM[16'h50EA] = 8'h00;
RAM[16'h50EB] = 8'h00;
RAM[16'h50EC] = 8'h00;
RAM[16'h50ED] = 8'h00;
RAM[16'h50EE] = 8'h00;
RAM[16'h50EF] = 8'h00;
RAM[16'h50F0] = 8'h00;
RAM[16'h50F1] = 8'h00;
RAM[16'h50F2] = 8'h00;
RAM[16'h50F3] = 8'h00;
RAM[16'h50F4] = 8'h00;
RAM[16'h50F5] = 8'h00;
RAM[16'h50F6] = 8'h00;
RAM[16'h50F7] = 8'h00;
RAM[16'h50F8] = 8'h00;
RAM[16'h50F9] = 8'h00;
RAM[16'h50FA] = 8'h00;
RAM[16'h50FB] = 8'h00;
RAM[16'h50FC] = 8'h00;
RAM[16'h50FD] = 8'h00;
RAM[16'h50FE] = 8'h00;
RAM[16'h50FF] = 8'h00;
RAM[16'h5100] = 8'h00;
RAM[16'h5101] = 8'h00;
RAM[16'h5102] = 8'h00;
RAM[16'h5103] = 8'h00;
RAM[16'h5104] = 8'h00;
RAM[16'h5105] = 8'h00;
RAM[16'h5106] = 8'h00;
RAM[16'h5107] = 8'h00;
RAM[16'h5108] = 8'h00;
RAM[16'h5109] = 8'h00;
RAM[16'h510A] = 8'h00;
RAM[16'h510B] = 8'h00;
RAM[16'h510C] = 8'h00;
RAM[16'h510D] = 8'h00;
RAM[16'h510E] = 8'h00;
RAM[16'h510F] = 8'h00;
RAM[16'h5110] = 8'h00;
RAM[16'h5111] = 8'h00;
RAM[16'h5112] = 8'h00;
RAM[16'h5113] = 8'h00;
RAM[16'h5114] = 8'h00;
RAM[16'h5115] = 8'h00;
RAM[16'h5116] = 8'h00;
RAM[16'h5117] = 8'h00;
RAM[16'h5118] = 8'h00;
RAM[16'h5119] = 8'h00;
RAM[16'h511A] = 8'h00;
RAM[16'h511B] = 8'h00;
RAM[16'h511C] = 8'h00;
RAM[16'h511D] = 8'h00;
RAM[16'h511E] = 8'h00;
RAM[16'h511F] = 8'h00;
RAM[16'h5120] = 8'h00;
RAM[16'h5121] = 8'h00;
RAM[16'h5122] = 8'h00;
RAM[16'h5123] = 8'h00;
RAM[16'h5124] = 8'h00;
RAM[16'h5125] = 8'h00;
RAM[16'h5126] = 8'h00;
RAM[16'h5127] = 8'h00;
RAM[16'h5128] = 8'h00;
RAM[16'h5129] = 8'h00;
RAM[16'h512A] = 8'h00;
RAM[16'h512B] = 8'h00;
RAM[16'h512C] = 8'h00;
RAM[16'h512D] = 8'h00;
RAM[16'h512E] = 8'h00;
RAM[16'h512F] = 8'h00;
RAM[16'h5130] = 8'h00;
RAM[16'h5131] = 8'h00;
RAM[16'h5132] = 8'h00;
RAM[16'h5133] = 8'h00;
RAM[16'h5134] = 8'h00;
RAM[16'h5135] = 8'h00;
RAM[16'h5136] = 8'h00;
RAM[16'h5137] = 8'h00;
RAM[16'h5138] = 8'h00;
RAM[16'h5139] = 8'h00;
RAM[16'h513A] = 8'h00;
RAM[16'h513B] = 8'h00;
RAM[16'h513C] = 8'h00;
RAM[16'h513D] = 8'h00;
RAM[16'h513E] = 8'h00;
RAM[16'h513F] = 8'h00;
RAM[16'h5140] = 8'h00;
RAM[16'h5141] = 8'h00;
RAM[16'h5142] = 8'h00;
RAM[16'h5143] = 8'h00;
RAM[16'h5144] = 8'h00;
RAM[16'h5145] = 8'h00;
RAM[16'h5146] = 8'h00;
RAM[16'h5147] = 8'h00;
RAM[16'h5148] = 8'h00;
RAM[16'h5149] = 8'h00;
RAM[16'h514A] = 8'h00;
RAM[16'h514B] = 8'h00;
RAM[16'h514C] = 8'h00;
RAM[16'h514D] = 8'h00;
RAM[16'h514E] = 8'h00;
RAM[16'h514F] = 8'h00;
RAM[16'h5150] = 8'h00;
RAM[16'h5151] = 8'h00;
RAM[16'h5152] = 8'h00;
RAM[16'h5153] = 8'h00;
RAM[16'h5154] = 8'h00;
RAM[16'h5155] = 8'h00;
RAM[16'h5156] = 8'h00;
RAM[16'h5157] = 8'h00;
RAM[16'h5158] = 8'h00;
RAM[16'h5159] = 8'h00;
RAM[16'h515A] = 8'h00;
RAM[16'h515B] = 8'h00;
RAM[16'h515C] = 8'h00;
RAM[16'h515D] = 8'h00;
RAM[16'h515E] = 8'h00;
RAM[16'h515F] = 8'h00;
RAM[16'h5160] = 8'h00;
RAM[16'h5161] = 8'h00;
RAM[16'h5162] = 8'h00;
RAM[16'h5163] = 8'h00;
RAM[16'h5164] = 8'h00;
RAM[16'h5165] = 8'h00;
RAM[16'h5166] = 8'h00;
RAM[16'h5167] = 8'h00;
RAM[16'h5168] = 8'h00;
RAM[16'h5169] = 8'h00;
RAM[16'h516A] = 8'h00;
RAM[16'h516B] = 8'h00;
RAM[16'h516C] = 8'h00;
RAM[16'h516D] = 8'h00;
RAM[16'h516E] = 8'h00;
RAM[16'h516F] = 8'h00;
RAM[16'h5170] = 8'h00;
RAM[16'h5171] = 8'h00;
RAM[16'h5172] = 8'h00;
RAM[16'h5173] = 8'h00;
RAM[16'h5174] = 8'h00;
RAM[16'h5175] = 8'h00;
RAM[16'h5176] = 8'h00;
RAM[16'h5177] = 8'h00;
RAM[16'h5178] = 8'h00;
RAM[16'h5179] = 8'h00;
RAM[16'h517A] = 8'h00;
RAM[16'h517B] = 8'h00;
RAM[16'h517C] = 8'h00;
RAM[16'h517D] = 8'h00;
RAM[16'h517E] = 8'h00;
RAM[16'h517F] = 8'h00;
RAM[16'h5180] = 8'h00;
RAM[16'h5181] = 8'h00;
RAM[16'h5182] = 8'h00;
RAM[16'h5183] = 8'h00;
RAM[16'h5184] = 8'h00;
RAM[16'h5185] = 8'h00;
RAM[16'h5186] = 8'h00;
RAM[16'h5187] = 8'h00;
RAM[16'h5188] = 8'h00;
RAM[16'h5189] = 8'h00;
RAM[16'h518A] = 8'h00;
RAM[16'h518B] = 8'h00;
RAM[16'h518C] = 8'h00;
RAM[16'h518D] = 8'h00;
RAM[16'h518E] = 8'h00;
RAM[16'h518F] = 8'h00;
RAM[16'h5190] = 8'h00;
RAM[16'h5191] = 8'h00;
RAM[16'h5192] = 8'h00;
RAM[16'h5193] = 8'h00;
RAM[16'h5194] = 8'h00;
RAM[16'h5195] = 8'h00;
RAM[16'h5196] = 8'h00;
RAM[16'h5197] = 8'h00;
RAM[16'h5198] = 8'h00;
RAM[16'h5199] = 8'h00;
RAM[16'h519A] = 8'h00;
RAM[16'h519B] = 8'h00;
RAM[16'h519C] = 8'h00;
RAM[16'h519D] = 8'h00;
RAM[16'h519E] = 8'h00;
RAM[16'h519F] = 8'h00;
RAM[16'h51A0] = 8'h00;
RAM[16'h51A1] = 8'h00;
RAM[16'h51A2] = 8'h00;
RAM[16'h51A3] = 8'h00;
RAM[16'h51A4] = 8'h00;
RAM[16'h51A5] = 8'h00;
RAM[16'h51A6] = 8'h00;
RAM[16'h51A7] = 8'h00;
RAM[16'h51A8] = 8'h00;
RAM[16'h51A9] = 8'h00;
RAM[16'h51AA] = 8'h00;
RAM[16'h51AB] = 8'h00;
RAM[16'h51AC] = 8'h00;
RAM[16'h51AD] = 8'h00;
RAM[16'h51AE] = 8'h00;
RAM[16'h51AF] = 8'h00;
RAM[16'h51B0] = 8'h00;
RAM[16'h51B1] = 8'h00;
RAM[16'h51B2] = 8'h00;
RAM[16'h51B3] = 8'h00;
RAM[16'h51B4] = 8'h00;
RAM[16'h51B5] = 8'h00;
RAM[16'h51B6] = 8'h00;
RAM[16'h51B7] = 8'h00;
RAM[16'h51B8] = 8'h00;
RAM[16'h51B9] = 8'h00;
RAM[16'h51BA] = 8'h00;
RAM[16'h51BB] = 8'h00;
RAM[16'h51BC] = 8'h00;
RAM[16'h51BD] = 8'h00;
RAM[16'h51BE] = 8'h00;
RAM[16'h51BF] = 8'h00;
RAM[16'h51C0] = 8'h00;
RAM[16'h51C1] = 8'h00;
RAM[16'h51C2] = 8'h00;
RAM[16'h51C3] = 8'h00;
RAM[16'h51C4] = 8'h00;
RAM[16'h51C5] = 8'h00;
RAM[16'h51C6] = 8'h00;
RAM[16'h51C7] = 8'h00;
RAM[16'h51C8] = 8'h00;
RAM[16'h51C9] = 8'h00;
RAM[16'h51CA] = 8'h00;
RAM[16'h51CB] = 8'h00;
RAM[16'h51CC] = 8'h00;
RAM[16'h51CD] = 8'h00;
RAM[16'h51CE] = 8'h00;
RAM[16'h51CF] = 8'h00;
RAM[16'h51D0] = 8'h00;
RAM[16'h51D1] = 8'h00;
RAM[16'h51D2] = 8'h00;
RAM[16'h51D3] = 8'h00;
RAM[16'h51D4] = 8'h00;
RAM[16'h51D5] = 8'h00;
RAM[16'h51D6] = 8'h00;
RAM[16'h51D7] = 8'h00;
RAM[16'h51D8] = 8'h00;
RAM[16'h51D9] = 8'h00;
RAM[16'h51DA] = 8'h00;
RAM[16'h51DB] = 8'h00;
RAM[16'h51DC] = 8'h00;
RAM[16'h51DD] = 8'h00;
RAM[16'h51DE] = 8'h00;
RAM[16'h51DF] = 8'h00;
RAM[16'h51E0] = 8'h00;
RAM[16'h51E1] = 8'h00;
RAM[16'h51E2] = 8'h00;
RAM[16'h51E3] = 8'h00;
RAM[16'h51E4] = 8'h00;
RAM[16'h51E5] = 8'h00;
RAM[16'h51E6] = 8'h00;
RAM[16'h51E7] = 8'h00;
RAM[16'h51E8] = 8'h00;
RAM[16'h51E9] = 8'h00;
RAM[16'h51EA] = 8'h00;
RAM[16'h51EB] = 8'h00;
RAM[16'h51EC] = 8'h00;
RAM[16'h51ED] = 8'h00;
RAM[16'h51EE] = 8'h00;
RAM[16'h51EF] = 8'h00;
RAM[16'h51F0] = 8'h00;
RAM[16'h51F1] = 8'h00;
RAM[16'h51F2] = 8'h00;
RAM[16'h51F3] = 8'h00;
RAM[16'h51F4] = 8'h00;
RAM[16'h51F5] = 8'h00;
RAM[16'h51F6] = 8'h00;
RAM[16'h51F7] = 8'h00;
RAM[16'h51F8] = 8'h00;
RAM[16'h51F9] = 8'h00;
RAM[16'h51FA] = 8'h00;
RAM[16'h51FB] = 8'h00;
RAM[16'h51FC] = 8'h00;
RAM[16'h51FD] = 8'h00;
RAM[16'h51FE] = 8'h00;
RAM[16'h51FF] = 8'h00;
RAM[16'h5200] = 8'h00;
RAM[16'h5201] = 8'h00;
RAM[16'h5202] = 8'h00;
RAM[16'h5203] = 8'h00;
RAM[16'h5204] = 8'h00;
RAM[16'h5205] = 8'h00;
RAM[16'h5206] = 8'h00;
RAM[16'h5207] = 8'h00;
RAM[16'h5208] = 8'h00;
RAM[16'h5209] = 8'h00;
RAM[16'h520A] = 8'h00;
RAM[16'h520B] = 8'h00;
RAM[16'h520C] = 8'h00;
RAM[16'h520D] = 8'h00;
RAM[16'h520E] = 8'h00;
RAM[16'h520F] = 8'h00;
RAM[16'h5210] = 8'h00;
RAM[16'h5211] = 8'h00;
RAM[16'h5212] = 8'h00;
RAM[16'h5213] = 8'h00;
RAM[16'h5214] = 8'h00;
RAM[16'h5215] = 8'h00;
RAM[16'h5216] = 8'h00;
RAM[16'h5217] = 8'h00;
RAM[16'h5218] = 8'h00;
RAM[16'h5219] = 8'h00;
RAM[16'h521A] = 8'h00;
RAM[16'h521B] = 8'h00;
RAM[16'h521C] = 8'h00;
RAM[16'h521D] = 8'h00;
RAM[16'h521E] = 8'h00;
RAM[16'h521F] = 8'h00;
RAM[16'h5220] = 8'h00;
RAM[16'h5221] = 8'h00;
RAM[16'h5222] = 8'h00;
RAM[16'h5223] = 8'h00;
RAM[16'h5224] = 8'h00;
RAM[16'h5225] = 8'h00;
RAM[16'h5226] = 8'h00;
RAM[16'h5227] = 8'h00;
RAM[16'h5228] = 8'h00;
RAM[16'h5229] = 8'h00;
RAM[16'h522A] = 8'h00;
RAM[16'h522B] = 8'h00;
RAM[16'h522C] = 8'h00;
RAM[16'h522D] = 8'h00;
RAM[16'h522E] = 8'h00;
RAM[16'h522F] = 8'h00;
RAM[16'h5230] = 8'h00;
RAM[16'h5231] = 8'h00;
RAM[16'h5232] = 8'h00;
RAM[16'h5233] = 8'h00;
RAM[16'h5234] = 8'h00;
RAM[16'h5235] = 8'h00;
RAM[16'h5236] = 8'h00;
RAM[16'h5237] = 8'h00;
RAM[16'h5238] = 8'h00;
RAM[16'h5239] = 8'h00;
RAM[16'h523A] = 8'h00;
RAM[16'h523B] = 8'h00;
RAM[16'h523C] = 8'h00;
RAM[16'h523D] = 8'h00;
RAM[16'h523E] = 8'h00;
RAM[16'h523F] = 8'h00;
RAM[16'h5240] = 8'h00;
RAM[16'h5241] = 8'h00;
RAM[16'h5242] = 8'h00;
RAM[16'h5243] = 8'h00;
RAM[16'h5244] = 8'h00;
RAM[16'h5245] = 8'h00;
RAM[16'h5246] = 8'h00;
RAM[16'h5247] = 8'h00;
RAM[16'h5248] = 8'h00;
RAM[16'h5249] = 8'h00;
RAM[16'h524A] = 8'h00;
RAM[16'h524B] = 8'h00;
RAM[16'h524C] = 8'h00;
RAM[16'h524D] = 8'h00;
RAM[16'h524E] = 8'h00;
RAM[16'h524F] = 8'h00;
RAM[16'h5250] = 8'h00;
RAM[16'h5251] = 8'h00;
RAM[16'h5252] = 8'h00;
RAM[16'h5253] = 8'h00;
RAM[16'h5254] = 8'h00;
RAM[16'h5255] = 8'h00;
RAM[16'h5256] = 8'h00;
RAM[16'h5257] = 8'h00;
RAM[16'h5258] = 8'h00;
RAM[16'h5259] = 8'h00;
RAM[16'h525A] = 8'h00;
RAM[16'h525B] = 8'h00;
RAM[16'h525C] = 8'h00;
RAM[16'h525D] = 8'h00;
RAM[16'h525E] = 8'h00;
RAM[16'h525F] = 8'h00;
RAM[16'h5260] = 8'h00;
RAM[16'h5261] = 8'h00;
RAM[16'h5262] = 8'h00;
RAM[16'h5263] = 8'h00;
RAM[16'h5264] = 8'h00;
RAM[16'h5265] = 8'h00;
RAM[16'h5266] = 8'h00;
RAM[16'h5267] = 8'h00;
RAM[16'h5268] = 8'h00;
RAM[16'h5269] = 8'h00;
RAM[16'h526A] = 8'h00;
RAM[16'h526B] = 8'h00;
RAM[16'h526C] = 8'h00;
RAM[16'h526D] = 8'h00;
RAM[16'h526E] = 8'h00;
RAM[16'h526F] = 8'h00;
RAM[16'h5270] = 8'h00;
RAM[16'h5271] = 8'h00;
RAM[16'h5272] = 8'h00;
RAM[16'h5273] = 8'h00;
RAM[16'h5274] = 8'h00;
RAM[16'h5275] = 8'h00;
RAM[16'h5276] = 8'h00;
RAM[16'h5277] = 8'h00;
RAM[16'h5278] = 8'h00;
RAM[16'h5279] = 8'h00;
RAM[16'h527A] = 8'h00;
RAM[16'h527B] = 8'h00;
RAM[16'h527C] = 8'h00;
RAM[16'h527D] = 8'h00;
RAM[16'h527E] = 8'h00;
RAM[16'h527F] = 8'h00;
RAM[16'h5280] = 8'h00;
RAM[16'h5281] = 8'h00;
RAM[16'h5282] = 8'h00;
RAM[16'h5283] = 8'h00;
RAM[16'h5284] = 8'h00;
RAM[16'h5285] = 8'h00;
RAM[16'h5286] = 8'h00;
RAM[16'h5287] = 8'h00;
RAM[16'h5288] = 8'h00;
RAM[16'h5289] = 8'h00;
RAM[16'h528A] = 8'h00;
RAM[16'h528B] = 8'h00;
RAM[16'h528C] = 8'h00;
RAM[16'h528D] = 8'h00;
RAM[16'h528E] = 8'h00;
RAM[16'h528F] = 8'h00;
RAM[16'h5290] = 8'h00;
RAM[16'h5291] = 8'h00;
RAM[16'h5292] = 8'h00;
RAM[16'h5293] = 8'h00;
RAM[16'h5294] = 8'h00;
RAM[16'h5295] = 8'h00;
RAM[16'h5296] = 8'h00;
RAM[16'h5297] = 8'h00;
RAM[16'h5298] = 8'h00;
RAM[16'h5299] = 8'h00;
RAM[16'h529A] = 8'h00;
RAM[16'h529B] = 8'h00;
RAM[16'h529C] = 8'h00;
RAM[16'h529D] = 8'h00;
RAM[16'h529E] = 8'h00;
RAM[16'h529F] = 8'h00;
RAM[16'h52A0] = 8'h00;
RAM[16'h52A1] = 8'h00;
RAM[16'h52A2] = 8'h00;
RAM[16'h52A3] = 8'h00;
RAM[16'h52A4] = 8'h00;
RAM[16'h52A5] = 8'h00;
RAM[16'h52A6] = 8'h00;
RAM[16'h52A7] = 8'h00;
RAM[16'h52A8] = 8'h00;
RAM[16'h52A9] = 8'h00;
RAM[16'h52AA] = 8'h00;
RAM[16'h52AB] = 8'h00;
RAM[16'h52AC] = 8'h00;
RAM[16'h52AD] = 8'h00;
RAM[16'h52AE] = 8'h00;
RAM[16'h52AF] = 8'h00;
RAM[16'h52B0] = 8'h00;
RAM[16'h52B1] = 8'h00;
RAM[16'h52B2] = 8'h00;
RAM[16'h52B3] = 8'h00;
RAM[16'h52B4] = 8'h00;
RAM[16'h52B5] = 8'h00;
RAM[16'h52B6] = 8'h00;
RAM[16'h52B7] = 8'h00;
RAM[16'h52B8] = 8'h00;
RAM[16'h52B9] = 8'h00;
RAM[16'h52BA] = 8'h00;
RAM[16'h52BB] = 8'h00;
RAM[16'h52BC] = 8'h00;
RAM[16'h52BD] = 8'h00;
RAM[16'h52BE] = 8'h00;
RAM[16'h52BF] = 8'h00;
RAM[16'h52C0] = 8'h00;
RAM[16'h52C1] = 8'h00;
RAM[16'h52C2] = 8'h00;
RAM[16'h52C3] = 8'h00;
RAM[16'h52C4] = 8'h00;
RAM[16'h52C5] = 8'h00;
RAM[16'h52C6] = 8'h00;
RAM[16'h52C7] = 8'h00;
RAM[16'h52C8] = 8'h00;
RAM[16'h52C9] = 8'h00;
RAM[16'h52CA] = 8'h00;
RAM[16'h52CB] = 8'h00;
RAM[16'h52CC] = 8'h00;
RAM[16'h52CD] = 8'h00;
RAM[16'h52CE] = 8'h00;
RAM[16'h52CF] = 8'h00;
RAM[16'h52D0] = 8'h00;
RAM[16'h52D1] = 8'h00;
RAM[16'h52D2] = 8'h00;
RAM[16'h52D3] = 8'h00;
RAM[16'h52D4] = 8'h00;
RAM[16'h52D5] = 8'h00;
RAM[16'h52D6] = 8'h00;
RAM[16'h52D7] = 8'h00;
RAM[16'h52D8] = 8'h00;
RAM[16'h52D9] = 8'h00;
RAM[16'h52DA] = 8'h00;
RAM[16'h52DB] = 8'h00;
RAM[16'h52DC] = 8'h00;
RAM[16'h52DD] = 8'h00;
RAM[16'h52DE] = 8'h00;
RAM[16'h52DF] = 8'h00;
RAM[16'h52E0] = 8'h00;
RAM[16'h52E1] = 8'h00;
RAM[16'h52E2] = 8'h00;
RAM[16'h52E3] = 8'h00;
RAM[16'h52E4] = 8'h00;
RAM[16'h52E5] = 8'h00;
RAM[16'h52E6] = 8'h00;
RAM[16'h52E7] = 8'h00;
RAM[16'h52E8] = 8'h00;
RAM[16'h52E9] = 8'h00;
RAM[16'h52EA] = 8'h00;
RAM[16'h52EB] = 8'h00;
RAM[16'h52EC] = 8'h00;
RAM[16'h52ED] = 8'h00;
RAM[16'h52EE] = 8'h00;
RAM[16'h52EF] = 8'h00;
RAM[16'h52F0] = 8'h00;
RAM[16'h52F1] = 8'h00;
RAM[16'h52F2] = 8'h00;
RAM[16'h52F3] = 8'h00;
RAM[16'h52F4] = 8'h00;
RAM[16'h52F5] = 8'h00;
RAM[16'h52F6] = 8'h00;
RAM[16'h52F7] = 8'h00;
RAM[16'h52F8] = 8'h00;
RAM[16'h52F9] = 8'h00;
RAM[16'h52FA] = 8'h00;
RAM[16'h52FB] = 8'h00;
RAM[16'h52FC] = 8'h00;
RAM[16'h52FD] = 8'h00;
RAM[16'h52FE] = 8'h00;
RAM[16'h52FF] = 8'h00;
RAM[16'h5300] = 8'h00;
RAM[16'h5301] = 8'h00;
RAM[16'h5302] = 8'h00;
RAM[16'h5303] = 8'h00;
RAM[16'h5304] = 8'h00;
RAM[16'h5305] = 8'h00;
RAM[16'h5306] = 8'h00;
RAM[16'h5307] = 8'h00;
RAM[16'h5308] = 8'h00;
RAM[16'h5309] = 8'h00;
RAM[16'h530A] = 8'h00;
RAM[16'h530B] = 8'h00;
RAM[16'h530C] = 8'h00;
RAM[16'h530D] = 8'h00;
RAM[16'h530E] = 8'h00;
RAM[16'h530F] = 8'h00;
RAM[16'h5310] = 8'h00;
RAM[16'h5311] = 8'h00;
RAM[16'h5312] = 8'h00;
RAM[16'h5313] = 8'h00;
RAM[16'h5314] = 8'h00;
RAM[16'h5315] = 8'h00;
RAM[16'h5316] = 8'h00;
RAM[16'h5317] = 8'h00;
RAM[16'h5318] = 8'h00;
RAM[16'h5319] = 8'h00;
RAM[16'h531A] = 8'h00;
RAM[16'h531B] = 8'h00;
RAM[16'h531C] = 8'h00;
RAM[16'h531D] = 8'h00;
RAM[16'h531E] = 8'h00;
RAM[16'h531F] = 8'h00;
RAM[16'h5320] = 8'h00;
RAM[16'h5321] = 8'h00;
RAM[16'h5322] = 8'h00;
RAM[16'h5323] = 8'h00;
RAM[16'h5324] = 8'h00;
RAM[16'h5325] = 8'h00;
RAM[16'h5326] = 8'h00;
RAM[16'h5327] = 8'h00;
RAM[16'h5328] = 8'h00;
RAM[16'h5329] = 8'h00;
RAM[16'h532A] = 8'h00;
RAM[16'h532B] = 8'h00;
RAM[16'h532C] = 8'h00;
RAM[16'h532D] = 8'h00;
RAM[16'h532E] = 8'h00;
RAM[16'h532F] = 8'h00;
RAM[16'h5330] = 8'h00;
RAM[16'h5331] = 8'h00;
RAM[16'h5332] = 8'h00;
RAM[16'h5333] = 8'h00;
RAM[16'h5334] = 8'h00;
RAM[16'h5335] = 8'h00;
RAM[16'h5336] = 8'h00;
RAM[16'h5337] = 8'h00;
RAM[16'h5338] = 8'h00;
RAM[16'h5339] = 8'h00;
RAM[16'h533A] = 8'h00;
RAM[16'h533B] = 8'h00;
RAM[16'h533C] = 8'h00;
RAM[16'h533D] = 8'h00;
RAM[16'h533E] = 8'h00;
RAM[16'h533F] = 8'h00;
RAM[16'h5340] = 8'h00;
RAM[16'h5341] = 8'h00;
RAM[16'h5342] = 8'h00;
RAM[16'h5343] = 8'h00;
RAM[16'h5344] = 8'h00;
RAM[16'h5345] = 8'h00;
RAM[16'h5346] = 8'h00;
RAM[16'h5347] = 8'h00;
RAM[16'h5348] = 8'h00;
RAM[16'h5349] = 8'h00;
RAM[16'h534A] = 8'h00;
RAM[16'h534B] = 8'h00;
RAM[16'h534C] = 8'h00;
RAM[16'h534D] = 8'h00;
RAM[16'h534E] = 8'h00;
RAM[16'h534F] = 8'h00;
RAM[16'h5350] = 8'h00;
RAM[16'h5351] = 8'h00;
RAM[16'h5352] = 8'h00;
RAM[16'h5353] = 8'h00;
RAM[16'h5354] = 8'h00;
RAM[16'h5355] = 8'h00;
RAM[16'h5356] = 8'h00;
RAM[16'h5357] = 8'h00;
RAM[16'h5358] = 8'h00;
RAM[16'h5359] = 8'h00;
RAM[16'h535A] = 8'h00;
RAM[16'h535B] = 8'h00;
RAM[16'h535C] = 8'h00;
RAM[16'h535D] = 8'h00;
RAM[16'h535E] = 8'h00;
RAM[16'h535F] = 8'h00;
RAM[16'h5360] = 8'h00;
RAM[16'h5361] = 8'h00;
RAM[16'h5362] = 8'h00;
RAM[16'h5363] = 8'h00;
RAM[16'h5364] = 8'h00;
RAM[16'h5365] = 8'h00;
RAM[16'h5366] = 8'h00;
RAM[16'h5367] = 8'h00;
RAM[16'h5368] = 8'h00;
RAM[16'h5369] = 8'h00;
RAM[16'h536A] = 8'h00;
RAM[16'h536B] = 8'h00;
RAM[16'h536C] = 8'h00;
RAM[16'h536D] = 8'h00;
RAM[16'h536E] = 8'h00;
RAM[16'h536F] = 8'h00;
RAM[16'h5370] = 8'h00;
RAM[16'h5371] = 8'h00;
RAM[16'h5372] = 8'h00;
RAM[16'h5373] = 8'h00;
RAM[16'h5374] = 8'h00;
RAM[16'h5375] = 8'h00;
RAM[16'h5376] = 8'h00;
RAM[16'h5377] = 8'h00;
RAM[16'h5378] = 8'h00;
RAM[16'h5379] = 8'h00;
RAM[16'h537A] = 8'h00;
RAM[16'h537B] = 8'h00;
RAM[16'h537C] = 8'h00;
RAM[16'h537D] = 8'h00;
RAM[16'h537E] = 8'h00;
RAM[16'h537F] = 8'h00;
RAM[16'h5380] = 8'h00;
RAM[16'h5381] = 8'h00;
RAM[16'h5382] = 8'h00;
RAM[16'h5383] = 8'h00;
RAM[16'h5384] = 8'h00;
RAM[16'h5385] = 8'h00;
RAM[16'h5386] = 8'h00;
RAM[16'h5387] = 8'h00;
RAM[16'h5388] = 8'h00;
RAM[16'h5389] = 8'h00;
RAM[16'h538A] = 8'h00;
RAM[16'h538B] = 8'h00;
RAM[16'h538C] = 8'h00;
RAM[16'h538D] = 8'h00;
RAM[16'h538E] = 8'h00;
RAM[16'h538F] = 8'h00;
RAM[16'h5390] = 8'h00;
RAM[16'h5391] = 8'h00;
RAM[16'h5392] = 8'h00;
RAM[16'h5393] = 8'h00;
RAM[16'h5394] = 8'h00;
RAM[16'h5395] = 8'h00;
RAM[16'h5396] = 8'h00;
RAM[16'h5397] = 8'h00;
RAM[16'h5398] = 8'h00;
RAM[16'h5399] = 8'h00;
RAM[16'h539A] = 8'h00;
RAM[16'h539B] = 8'h00;
RAM[16'h539C] = 8'h00;
RAM[16'h539D] = 8'h00;
RAM[16'h539E] = 8'h00;
RAM[16'h539F] = 8'h00;
RAM[16'h53A0] = 8'h00;
RAM[16'h53A1] = 8'h00;
RAM[16'h53A2] = 8'h00;
RAM[16'h53A3] = 8'h00;
RAM[16'h53A4] = 8'h00;
RAM[16'h53A5] = 8'h00;
RAM[16'h53A6] = 8'h00;
RAM[16'h53A7] = 8'h00;
RAM[16'h53A8] = 8'h00;
RAM[16'h53A9] = 8'h00;
RAM[16'h53AA] = 8'h00;
RAM[16'h53AB] = 8'h00;
RAM[16'h53AC] = 8'h00;
RAM[16'h53AD] = 8'h00;
RAM[16'h53AE] = 8'h00;
RAM[16'h53AF] = 8'h00;
RAM[16'h53B0] = 8'h00;
RAM[16'h53B1] = 8'h00;
RAM[16'h53B2] = 8'h00;
RAM[16'h53B3] = 8'h00;
RAM[16'h53B4] = 8'h00;
RAM[16'h53B5] = 8'h00;
RAM[16'h53B6] = 8'h00;
RAM[16'h53B7] = 8'h00;
RAM[16'h53B8] = 8'h00;
RAM[16'h53B9] = 8'h00;
RAM[16'h53BA] = 8'h00;
RAM[16'h53BB] = 8'h00;
RAM[16'h53BC] = 8'h00;
RAM[16'h53BD] = 8'h00;
RAM[16'h53BE] = 8'h00;
RAM[16'h53BF] = 8'h00;
RAM[16'h53C0] = 8'h00;
RAM[16'h53C1] = 8'h00;
RAM[16'h53C2] = 8'h00;
RAM[16'h53C3] = 8'h00;
RAM[16'h53C4] = 8'h00;
RAM[16'h53C5] = 8'h00;
RAM[16'h53C6] = 8'h00;
RAM[16'h53C7] = 8'h00;
RAM[16'h53C8] = 8'h00;
RAM[16'h53C9] = 8'h00;
RAM[16'h53CA] = 8'h00;
RAM[16'h53CB] = 8'h00;
RAM[16'h53CC] = 8'h00;
RAM[16'h53CD] = 8'h00;
RAM[16'h53CE] = 8'h00;
RAM[16'h53CF] = 8'h00;
RAM[16'h53D0] = 8'h00;
RAM[16'h53D1] = 8'h00;
RAM[16'h53D2] = 8'h00;
RAM[16'h53D3] = 8'h00;
RAM[16'h53D4] = 8'h00;
RAM[16'h53D5] = 8'h00;
RAM[16'h53D6] = 8'h00;
RAM[16'h53D7] = 8'h00;
RAM[16'h53D8] = 8'h00;
RAM[16'h53D9] = 8'h00;
RAM[16'h53DA] = 8'h00;
RAM[16'h53DB] = 8'h00;
RAM[16'h53DC] = 8'h00;
RAM[16'h53DD] = 8'h00;
RAM[16'h53DE] = 8'h00;
RAM[16'h53DF] = 8'h00;
RAM[16'h53E0] = 8'h00;
RAM[16'h53E1] = 8'h00;
RAM[16'h53E2] = 8'h00;
RAM[16'h53E3] = 8'h00;
RAM[16'h53E4] = 8'h00;
RAM[16'h53E5] = 8'h00;
RAM[16'h53E6] = 8'h00;
RAM[16'h53E7] = 8'h00;
RAM[16'h53E8] = 8'h00;
RAM[16'h53E9] = 8'h00;
RAM[16'h53EA] = 8'h00;
RAM[16'h53EB] = 8'h00;
RAM[16'h53EC] = 8'h00;
RAM[16'h53ED] = 8'h00;
RAM[16'h53EE] = 8'h00;
RAM[16'h53EF] = 8'h00;
RAM[16'h53F0] = 8'h00;
RAM[16'h53F1] = 8'h00;
RAM[16'h53F2] = 8'h00;
RAM[16'h53F3] = 8'h00;
RAM[16'h53F4] = 8'h00;
RAM[16'h53F5] = 8'h00;
RAM[16'h53F6] = 8'h00;
RAM[16'h53F7] = 8'h00;
RAM[16'h53F8] = 8'h00;
RAM[16'h53F9] = 8'h00;
RAM[16'h53FA] = 8'h00;
RAM[16'h53FB] = 8'h00;
RAM[16'h53FC] = 8'h00;
RAM[16'h53FD] = 8'h00;
RAM[16'h53FE] = 8'h00;
RAM[16'h53FF] = 8'h00;
RAM[16'h5400] = 8'h00;
RAM[16'h5401] = 8'h00;
RAM[16'h5402] = 8'h00;
RAM[16'h5403] = 8'h00;
RAM[16'h5404] = 8'h00;
RAM[16'h5405] = 8'h00;
RAM[16'h5406] = 8'h00;
RAM[16'h5407] = 8'h00;
RAM[16'h5408] = 8'h00;
RAM[16'h5409] = 8'h00;
RAM[16'h540A] = 8'h00;
RAM[16'h540B] = 8'h00;
RAM[16'h540C] = 8'h00;
RAM[16'h540D] = 8'h00;
RAM[16'h540E] = 8'h00;
RAM[16'h540F] = 8'h00;
RAM[16'h5410] = 8'h00;
RAM[16'h5411] = 8'h00;
RAM[16'h5412] = 8'h00;
RAM[16'h5413] = 8'h00;
RAM[16'h5414] = 8'h00;
RAM[16'h5415] = 8'h00;
RAM[16'h5416] = 8'h00;
RAM[16'h5417] = 8'h00;
RAM[16'h5418] = 8'h00;
RAM[16'h5419] = 8'h00;
RAM[16'h541A] = 8'h00;
RAM[16'h541B] = 8'h00;
RAM[16'h541C] = 8'h00;
RAM[16'h541D] = 8'h00;
RAM[16'h541E] = 8'h00;
RAM[16'h541F] = 8'h00;
RAM[16'h5420] = 8'h00;
RAM[16'h5421] = 8'h00;
RAM[16'h5422] = 8'h00;
RAM[16'h5423] = 8'h00;
RAM[16'h5424] = 8'h00;
RAM[16'h5425] = 8'h00;
RAM[16'h5426] = 8'h00;
RAM[16'h5427] = 8'h00;
RAM[16'h5428] = 8'h00;
RAM[16'h5429] = 8'h00;
RAM[16'h542A] = 8'h00;
RAM[16'h542B] = 8'h00;
RAM[16'h542C] = 8'h00;
RAM[16'h542D] = 8'h00;
RAM[16'h542E] = 8'h00;
RAM[16'h542F] = 8'h00;
RAM[16'h5430] = 8'h00;
RAM[16'h5431] = 8'h00;
RAM[16'h5432] = 8'h00;
RAM[16'h5433] = 8'h00;
RAM[16'h5434] = 8'h00;
RAM[16'h5435] = 8'h00;
RAM[16'h5436] = 8'h00;
RAM[16'h5437] = 8'h00;
RAM[16'h5438] = 8'h00;
RAM[16'h5439] = 8'h00;
RAM[16'h543A] = 8'h00;
RAM[16'h543B] = 8'h00;
RAM[16'h543C] = 8'h00;
RAM[16'h543D] = 8'h00;
RAM[16'h543E] = 8'h00;
RAM[16'h543F] = 8'h00;
RAM[16'h5440] = 8'h00;
RAM[16'h5441] = 8'h00;
RAM[16'h5442] = 8'h00;
RAM[16'h5443] = 8'h00;
RAM[16'h5444] = 8'h00;
RAM[16'h5445] = 8'h00;
RAM[16'h5446] = 8'h00;
RAM[16'h5447] = 8'h00;
RAM[16'h5448] = 8'h00;
RAM[16'h5449] = 8'h00;
RAM[16'h544A] = 8'h00;
RAM[16'h544B] = 8'h00;
RAM[16'h544C] = 8'h00;
RAM[16'h544D] = 8'h00;
RAM[16'h544E] = 8'h00;
RAM[16'h544F] = 8'h00;
RAM[16'h5450] = 8'h00;
RAM[16'h5451] = 8'h00;
RAM[16'h5452] = 8'h00;
RAM[16'h5453] = 8'h00;
RAM[16'h5454] = 8'h00;
RAM[16'h5455] = 8'h00;
RAM[16'h5456] = 8'h00;
RAM[16'h5457] = 8'h00;
RAM[16'h5458] = 8'h00;
RAM[16'h5459] = 8'h00;
RAM[16'h545A] = 8'h00;
RAM[16'h545B] = 8'h00;
RAM[16'h545C] = 8'h00;
RAM[16'h545D] = 8'h00;
RAM[16'h545E] = 8'h00;
RAM[16'h545F] = 8'h00;
RAM[16'h5460] = 8'h00;
RAM[16'h5461] = 8'h00;
RAM[16'h5462] = 8'h00;
RAM[16'h5463] = 8'h00;
RAM[16'h5464] = 8'h00;
RAM[16'h5465] = 8'h00;
RAM[16'h5466] = 8'h00;
RAM[16'h5467] = 8'h00;
RAM[16'h5468] = 8'h00;
RAM[16'h5469] = 8'h00;
RAM[16'h546A] = 8'h00;
RAM[16'h546B] = 8'h00;
RAM[16'h546C] = 8'h00;
RAM[16'h546D] = 8'h00;
RAM[16'h546E] = 8'h00;
RAM[16'h546F] = 8'h00;
RAM[16'h5470] = 8'h00;
RAM[16'h5471] = 8'h00;
RAM[16'h5472] = 8'h00;
RAM[16'h5473] = 8'h00;
RAM[16'h5474] = 8'h00;
RAM[16'h5475] = 8'h00;
RAM[16'h5476] = 8'h00;
RAM[16'h5477] = 8'h00;
RAM[16'h5478] = 8'h00;
RAM[16'h5479] = 8'h00;
RAM[16'h547A] = 8'h00;
RAM[16'h547B] = 8'h00;
RAM[16'h547C] = 8'h00;
RAM[16'h547D] = 8'h00;
RAM[16'h547E] = 8'h00;
RAM[16'h547F] = 8'h00;
RAM[16'h5480] = 8'h00;
RAM[16'h5481] = 8'h00;
RAM[16'h5482] = 8'h00;
RAM[16'h5483] = 8'h00;
RAM[16'h5484] = 8'h00;
RAM[16'h5485] = 8'h00;
RAM[16'h5486] = 8'h00;
RAM[16'h5487] = 8'h00;
RAM[16'h5488] = 8'h00;
RAM[16'h5489] = 8'h00;
RAM[16'h548A] = 8'h00;
RAM[16'h548B] = 8'h00;
RAM[16'h548C] = 8'h00;
RAM[16'h548D] = 8'h00;
RAM[16'h548E] = 8'h00;
RAM[16'h548F] = 8'h00;
RAM[16'h5490] = 8'h00;
RAM[16'h5491] = 8'h00;
RAM[16'h5492] = 8'h00;
RAM[16'h5493] = 8'h00;
RAM[16'h5494] = 8'h00;
RAM[16'h5495] = 8'h00;
RAM[16'h5496] = 8'h00;
RAM[16'h5497] = 8'h00;
RAM[16'h5498] = 8'h00;
RAM[16'h5499] = 8'h00;
RAM[16'h549A] = 8'h00;
RAM[16'h549B] = 8'h00;
RAM[16'h549C] = 8'h00;
RAM[16'h549D] = 8'h00;
RAM[16'h549E] = 8'h00;
RAM[16'h549F] = 8'h00;
RAM[16'h54A0] = 8'h00;
RAM[16'h54A1] = 8'h00;
RAM[16'h54A2] = 8'h00;
RAM[16'h54A3] = 8'h00;
RAM[16'h54A4] = 8'h00;
RAM[16'h54A5] = 8'h00;
RAM[16'h54A6] = 8'h00;
RAM[16'h54A7] = 8'h00;
RAM[16'h54A8] = 8'h00;
RAM[16'h54A9] = 8'h00;
RAM[16'h54AA] = 8'h00;
RAM[16'h54AB] = 8'h00;
RAM[16'h54AC] = 8'h00;
RAM[16'h54AD] = 8'h00;
RAM[16'h54AE] = 8'h00;
RAM[16'h54AF] = 8'h00;
RAM[16'h54B0] = 8'h00;
RAM[16'h54B1] = 8'h00;
RAM[16'h54B2] = 8'h00;
RAM[16'h54B3] = 8'h00;
RAM[16'h54B4] = 8'h00;
RAM[16'h54B5] = 8'h00;
RAM[16'h54B6] = 8'h00;
RAM[16'h54B7] = 8'h00;
RAM[16'h54B8] = 8'h00;
RAM[16'h54B9] = 8'h00;
RAM[16'h54BA] = 8'h00;
RAM[16'h54BB] = 8'h00;
RAM[16'h54BC] = 8'h00;
RAM[16'h54BD] = 8'h00;
RAM[16'h54BE] = 8'h00;
RAM[16'h54BF] = 8'h00;
RAM[16'h54C0] = 8'h00;
RAM[16'h54C1] = 8'h00;
RAM[16'h54C2] = 8'h00;
RAM[16'h54C3] = 8'h00;
RAM[16'h54C4] = 8'h00;
RAM[16'h54C5] = 8'h00;
RAM[16'h54C6] = 8'h00;
RAM[16'h54C7] = 8'h00;
RAM[16'h54C8] = 8'h00;
RAM[16'h54C9] = 8'h00;
RAM[16'h54CA] = 8'h00;
RAM[16'h54CB] = 8'h00;
RAM[16'h54CC] = 8'h00;
RAM[16'h54CD] = 8'h00;
RAM[16'h54CE] = 8'h00;
RAM[16'h54CF] = 8'h00;
RAM[16'h54D0] = 8'h00;
RAM[16'h54D1] = 8'h00;
RAM[16'h54D2] = 8'h00;
RAM[16'h54D3] = 8'h00;
RAM[16'h54D4] = 8'h00;
RAM[16'h54D5] = 8'h00;
RAM[16'h54D6] = 8'h00;
RAM[16'h54D7] = 8'h00;
RAM[16'h54D8] = 8'h00;
RAM[16'h54D9] = 8'h00;
RAM[16'h54DA] = 8'h00;
RAM[16'h54DB] = 8'h00;
RAM[16'h54DC] = 8'h00;
RAM[16'h54DD] = 8'h00;
RAM[16'h54DE] = 8'h00;
RAM[16'h54DF] = 8'h00;
RAM[16'h54E0] = 8'h00;
RAM[16'h54E1] = 8'h00;
RAM[16'h54E2] = 8'h00;
RAM[16'h54E3] = 8'h00;
RAM[16'h54E4] = 8'h00;
RAM[16'h54E5] = 8'h00;
RAM[16'h54E6] = 8'h00;
RAM[16'h54E7] = 8'h00;
RAM[16'h54E8] = 8'h00;
RAM[16'h54E9] = 8'h00;
RAM[16'h54EA] = 8'h00;
RAM[16'h54EB] = 8'h00;
RAM[16'h54EC] = 8'h00;
RAM[16'h54ED] = 8'h00;
RAM[16'h54EE] = 8'h00;
RAM[16'h54EF] = 8'h00;
RAM[16'h54F0] = 8'h00;
RAM[16'h54F1] = 8'h00;
RAM[16'h54F2] = 8'h00;
RAM[16'h54F3] = 8'h00;
RAM[16'h54F4] = 8'h00;
RAM[16'h54F5] = 8'h00;
RAM[16'h54F6] = 8'h00;
RAM[16'h54F7] = 8'h00;
RAM[16'h54F8] = 8'h00;
RAM[16'h54F9] = 8'h00;
RAM[16'h54FA] = 8'h00;
RAM[16'h54FB] = 8'h00;
RAM[16'h54FC] = 8'h00;
RAM[16'h54FD] = 8'h00;
RAM[16'h54FE] = 8'h00;
RAM[16'h54FF] = 8'h00;
RAM[16'h5500] = 8'h00;
RAM[16'h5501] = 8'h00;
RAM[16'h5502] = 8'h00;
RAM[16'h5503] = 8'h00;
RAM[16'h5504] = 8'h00;
RAM[16'h5505] = 8'h00;
RAM[16'h5506] = 8'h00;
RAM[16'h5507] = 8'h00;
RAM[16'h5508] = 8'h00;
RAM[16'h5509] = 8'h00;
RAM[16'h550A] = 8'h00;
RAM[16'h550B] = 8'h00;
RAM[16'h550C] = 8'h00;
RAM[16'h550D] = 8'h00;
RAM[16'h550E] = 8'h00;
RAM[16'h550F] = 8'h00;
RAM[16'h5510] = 8'h00;
RAM[16'h5511] = 8'h00;
RAM[16'h5512] = 8'h00;
RAM[16'h5513] = 8'h00;
RAM[16'h5514] = 8'h00;
RAM[16'h5515] = 8'h00;
RAM[16'h5516] = 8'h00;
RAM[16'h5517] = 8'h00;
RAM[16'h5518] = 8'h00;
RAM[16'h5519] = 8'h00;
RAM[16'h551A] = 8'h00;
RAM[16'h551B] = 8'h00;
RAM[16'h551C] = 8'h00;
RAM[16'h551D] = 8'h00;
RAM[16'h551E] = 8'h00;
RAM[16'h551F] = 8'h00;
RAM[16'h5520] = 8'h00;
RAM[16'h5521] = 8'h00;
RAM[16'h5522] = 8'h00;
RAM[16'h5523] = 8'h00;
RAM[16'h5524] = 8'h00;
RAM[16'h5525] = 8'h00;
RAM[16'h5526] = 8'h00;
RAM[16'h5527] = 8'h00;
RAM[16'h5528] = 8'h00;
RAM[16'h5529] = 8'h00;
RAM[16'h552A] = 8'h00;
RAM[16'h552B] = 8'h00;
RAM[16'h552C] = 8'h00;
RAM[16'h552D] = 8'h00;
RAM[16'h552E] = 8'h00;
RAM[16'h552F] = 8'h00;
RAM[16'h5530] = 8'h00;
RAM[16'h5531] = 8'h00;
RAM[16'h5532] = 8'h00;
RAM[16'h5533] = 8'h00;
RAM[16'h5534] = 8'h00;
RAM[16'h5535] = 8'h00;
RAM[16'h5536] = 8'h00;
RAM[16'h5537] = 8'h00;
RAM[16'h5538] = 8'h00;
RAM[16'h5539] = 8'h00;
RAM[16'h553A] = 8'h00;
RAM[16'h553B] = 8'h00;
RAM[16'h553C] = 8'h00;
RAM[16'h553D] = 8'h00;
RAM[16'h553E] = 8'h00;
RAM[16'h553F] = 8'h00;
RAM[16'h5540] = 8'h00;
RAM[16'h5541] = 8'h00;
RAM[16'h5542] = 8'h00;
RAM[16'h5543] = 8'h00;
RAM[16'h5544] = 8'h00;
RAM[16'h5545] = 8'h00;
RAM[16'h5546] = 8'h00;
RAM[16'h5547] = 8'h00;
RAM[16'h5548] = 8'h00;
RAM[16'h5549] = 8'h00;
RAM[16'h554A] = 8'h00;
RAM[16'h554B] = 8'h00;
RAM[16'h554C] = 8'h00;
RAM[16'h554D] = 8'h00;
RAM[16'h554E] = 8'h00;
RAM[16'h554F] = 8'h00;
RAM[16'h5550] = 8'h00;
RAM[16'h5551] = 8'h00;
RAM[16'h5552] = 8'h00;
RAM[16'h5553] = 8'h00;
RAM[16'h5554] = 8'h00;
RAM[16'h5555] = 8'h00;
RAM[16'h5556] = 8'h00;
RAM[16'h5557] = 8'h00;
RAM[16'h5558] = 8'h00;
RAM[16'h5559] = 8'h00;
RAM[16'h555A] = 8'h00;
RAM[16'h555B] = 8'h00;
RAM[16'h555C] = 8'h00;
RAM[16'h555D] = 8'h00;
RAM[16'h555E] = 8'h00;
RAM[16'h555F] = 8'h00;
RAM[16'h5560] = 8'h00;
RAM[16'h5561] = 8'h00;
RAM[16'h5562] = 8'h00;
RAM[16'h5563] = 8'h00;
RAM[16'h5564] = 8'h00;
RAM[16'h5565] = 8'h00;
RAM[16'h5566] = 8'h00;
RAM[16'h5567] = 8'h00;
RAM[16'h5568] = 8'h00;
RAM[16'h5569] = 8'h00;
RAM[16'h556A] = 8'h00;
RAM[16'h556B] = 8'h00;
RAM[16'h556C] = 8'h00;
RAM[16'h556D] = 8'h00;
RAM[16'h556E] = 8'h00;
RAM[16'h556F] = 8'h00;
RAM[16'h5570] = 8'h00;
RAM[16'h5571] = 8'h00;
RAM[16'h5572] = 8'h00;
RAM[16'h5573] = 8'h00;
RAM[16'h5574] = 8'h00;
RAM[16'h5575] = 8'h00;
RAM[16'h5576] = 8'h00;
RAM[16'h5577] = 8'h00;
RAM[16'h5578] = 8'h00;
RAM[16'h5579] = 8'h00;
RAM[16'h557A] = 8'h00;
RAM[16'h557B] = 8'h00;
RAM[16'h557C] = 8'h00;
RAM[16'h557D] = 8'h00;
RAM[16'h557E] = 8'h00;
RAM[16'h557F] = 8'h00;
RAM[16'h5580] = 8'h00;
RAM[16'h5581] = 8'h00;
RAM[16'h5582] = 8'h00;
RAM[16'h5583] = 8'h00;
RAM[16'h5584] = 8'h00;
RAM[16'h5585] = 8'h00;
RAM[16'h5586] = 8'h00;
RAM[16'h5587] = 8'h00;
RAM[16'h5588] = 8'h00;
RAM[16'h5589] = 8'h00;
RAM[16'h558A] = 8'h00;
RAM[16'h558B] = 8'h00;
RAM[16'h558C] = 8'h00;
RAM[16'h558D] = 8'h00;
RAM[16'h558E] = 8'h00;
RAM[16'h558F] = 8'h00;
RAM[16'h5590] = 8'h00;
RAM[16'h5591] = 8'h00;
RAM[16'h5592] = 8'h00;
RAM[16'h5593] = 8'h00;
RAM[16'h5594] = 8'h00;
RAM[16'h5595] = 8'h00;
RAM[16'h5596] = 8'h00;
RAM[16'h5597] = 8'h00;
RAM[16'h5598] = 8'h00;
RAM[16'h5599] = 8'h00;
RAM[16'h559A] = 8'h00;
RAM[16'h559B] = 8'h00;
RAM[16'h559C] = 8'h00;
RAM[16'h559D] = 8'h00;
RAM[16'h559E] = 8'h00;
RAM[16'h559F] = 8'h00;
RAM[16'h55A0] = 8'h00;
RAM[16'h55A1] = 8'h00;
RAM[16'h55A2] = 8'h00;
RAM[16'h55A3] = 8'h00;
RAM[16'h55A4] = 8'h00;
RAM[16'h55A5] = 8'h00;
RAM[16'h55A6] = 8'h00;
RAM[16'h55A7] = 8'h00;
RAM[16'h55A8] = 8'h00;
RAM[16'h55A9] = 8'h00;
RAM[16'h55AA] = 8'h00;
RAM[16'h55AB] = 8'h00;
RAM[16'h55AC] = 8'h00;
RAM[16'h55AD] = 8'h00;
RAM[16'h55AE] = 8'h00;
RAM[16'h55AF] = 8'h00;
RAM[16'h55B0] = 8'h00;
RAM[16'h55B1] = 8'h00;
RAM[16'h55B2] = 8'h00;
RAM[16'h55B3] = 8'h00;
RAM[16'h55B4] = 8'h00;
RAM[16'h55B5] = 8'h00;
RAM[16'h55B6] = 8'h00;
RAM[16'h55B7] = 8'h00;
RAM[16'h55B8] = 8'h00;
RAM[16'h55B9] = 8'h00;
RAM[16'h55BA] = 8'h00;
RAM[16'h55BB] = 8'h00;
RAM[16'h55BC] = 8'h00;
RAM[16'h55BD] = 8'h00;
RAM[16'h55BE] = 8'h00;
RAM[16'h55BF] = 8'h00;
RAM[16'h55C0] = 8'h00;
RAM[16'h55C1] = 8'h00;
RAM[16'h55C2] = 8'h00;
RAM[16'h55C3] = 8'h00;
RAM[16'h55C4] = 8'h00;
RAM[16'h55C5] = 8'h00;
RAM[16'h55C6] = 8'h00;
RAM[16'h55C7] = 8'h00;
RAM[16'h55C8] = 8'h00;
RAM[16'h55C9] = 8'h00;
RAM[16'h55CA] = 8'h00;
RAM[16'h55CB] = 8'h00;
RAM[16'h55CC] = 8'h00;
RAM[16'h55CD] = 8'h00;
RAM[16'h55CE] = 8'h00;
RAM[16'h55CF] = 8'h00;
RAM[16'h55D0] = 8'h00;
RAM[16'h55D1] = 8'h00;
RAM[16'h55D2] = 8'h00;
RAM[16'h55D3] = 8'h00;
RAM[16'h55D4] = 8'h00;
RAM[16'h55D5] = 8'h00;
RAM[16'h55D6] = 8'h00;
RAM[16'h55D7] = 8'h00;
RAM[16'h55D8] = 8'h00;
RAM[16'h55D9] = 8'h00;
RAM[16'h55DA] = 8'h00;
RAM[16'h55DB] = 8'h00;
RAM[16'h55DC] = 8'h00;
RAM[16'h55DD] = 8'h00;
RAM[16'h55DE] = 8'h00;
RAM[16'h55DF] = 8'h00;
RAM[16'h55E0] = 8'h00;
RAM[16'h55E1] = 8'h00;
RAM[16'h55E2] = 8'h00;
RAM[16'h55E3] = 8'h00;
RAM[16'h55E4] = 8'h00;
RAM[16'h55E5] = 8'h00;
RAM[16'h55E6] = 8'h00;
RAM[16'h55E7] = 8'h00;
RAM[16'h55E8] = 8'h00;
RAM[16'h55E9] = 8'h00;
RAM[16'h55EA] = 8'h00;
RAM[16'h55EB] = 8'h00;
RAM[16'h55EC] = 8'h00;
RAM[16'h55ED] = 8'h00;
RAM[16'h55EE] = 8'h00;
RAM[16'h55EF] = 8'h00;
RAM[16'h55F0] = 8'h00;
RAM[16'h55F1] = 8'h00;
RAM[16'h55F2] = 8'h00;
RAM[16'h55F3] = 8'h00;
RAM[16'h55F4] = 8'h00;
RAM[16'h55F5] = 8'h00;
RAM[16'h55F6] = 8'h00;
RAM[16'h55F7] = 8'h00;
RAM[16'h55F8] = 8'h00;
RAM[16'h55F9] = 8'h00;
RAM[16'h55FA] = 8'h00;
RAM[16'h55FB] = 8'h00;
RAM[16'h55FC] = 8'h00;
RAM[16'h55FD] = 8'h00;
RAM[16'h55FE] = 8'h00;
RAM[16'h55FF] = 8'h00;
RAM[16'h5600] = 8'h00;
RAM[16'h5601] = 8'h00;
RAM[16'h5602] = 8'h00;
RAM[16'h5603] = 8'h00;
RAM[16'h5604] = 8'h00;
RAM[16'h5605] = 8'h00;
RAM[16'h5606] = 8'h00;
RAM[16'h5607] = 8'h00;
RAM[16'h5608] = 8'h00;
RAM[16'h5609] = 8'h00;
RAM[16'h560A] = 8'h00;
RAM[16'h560B] = 8'h00;
RAM[16'h560C] = 8'h00;
RAM[16'h560D] = 8'h00;
RAM[16'h560E] = 8'h00;
RAM[16'h560F] = 8'h00;
RAM[16'h5610] = 8'h00;
RAM[16'h5611] = 8'h00;
RAM[16'h5612] = 8'h00;
RAM[16'h5613] = 8'h00;
RAM[16'h5614] = 8'h00;
RAM[16'h5615] = 8'h00;
RAM[16'h5616] = 8'h00;
RAM[16'h5617] = 8'h00;
RAM[16'h5618] = 8'h00;
RAM[16'h5619] = 8'h00;
RAM[16'h561A] = 8'h00;
RAM[16'h561B] = 8'h00;
RAM[16'h561C] = 8'h00;
RAM[16'h561D] = 8'h00;
RAM[16'h561E] = 8'h00;
RAM[16'h561F] = 8'h00;
RAM[16'h5620] = 8'h00;
RAM[16'h5621] = 8'h00;
RAM[16'h5622] = 8'h00;
RAM[16'h5623] = 8'h00;
RAM[16'h5624] = 8'h00;
RAM[16'h5625] = 8'h00;
RAM[16'h5626] = 8'h00;
RAM[16'h5627] = 8'h00;
RAM[16'h5628] = 8'h00;
RAM[16'h5629] = 8'h00;
RAM[16'h562A] = 8'h00;
RAM[16'h562B] = 8'h00;
RAM[16'h562C] = 8'h00;
RAM[16'h562D] = 8'h00;
RAM[16'h562E] = 8'h00;
RAM[16'h562F] = 8'h00;
RAM[16'h5630] = 8'h00;
RAM[16'h5631] = 8'h00;
RAM[16'h5632] = 8'h00;
RAM[16'h5633] = 8'h00;
RAM[16'h5634] = 8'h00;
RAM[16'h5635] = 8'h00;
RAM[16'h5636] = 8'h00;
RAM[16'h5637] = 8'h00;
RAM[16'h5638] = 8'h00;
RAM[16'h5639] = 8'h00;
RAM[16'h563A] = 8'h00;
RAM[16'h563B] = 8'h00;
RAM[16'h563C] = 8'h00;
RAM[16'h563D] = 8'h00;
RAM[16'h563E] = 8'h00;
RAM[16'h563F] = 8'h00;
RAM[16'h5640] = 8'h00;
RAM[16'h5641] = 8'h00;
RAM[16'h5642] = 8'h00;
RAM[16'h5643] = 8'h00;
RAM[16'h5644] = 8'h00;
RAM[16'h5645] = 8'h00;
RAM[16'h5646] = 8'h00;
RAM[16'h5647] = 8'h00;
RAM[16'h5648] = 8'h00;
RAM[16'h5649] = 8'h00;
RAM[16'h564A] = 8'h00;
RAM[16'h564B] = 8'h00;
RAM[16'h564C] = 8'h00;
RAM[16'h564D] = 8'h00;
RAM[16'h564E] = 8'h00;
RAM[16'h564F] = 8'h00;
RAM[16'h5650] = 8'h00;
RAM[16'h5651] = 8'h00;
RAM[16'h5652] = 8'h00;
RAM[16'h5653] = 8'h00;
RAM[16'h5654] = 8'h00;
RAM[16'h5655] = 8'h00;
RAM[16'h5656] = 8'h00;
RAM[16'h5657] = 8'h00;
RAM[16'h5658] = 8'h00;
RAM[16'h5659] = 8'h00;
RAM[16'h565A] = 8'h00;
RAM[16'h565B] = 8'h00;
RAM[16'h565C] = 8'h00;
RAM[16'h565D] = 8'h00;
RAM[16'h565E] = 8'h00;
RAM[16'h565F] = 8'h00;
RAM[16'h5660] = 8'h00;
RAM[16'h5661] = 8'h00;
RAM[16'h5662] = 8'h00;
RAM[16'h5663] = 8'h00;
RAM[16'h5664] = 8'h00;
RAM[16'h5665] = 8'h00;
RAM[16'h5666] = 8'h00;
RAM[16'h5667] = 8'h00;
RAM[16'h5668] = 8'h00;
RAM[16'h5669] = 8'h00;
RAM[16'h566A] = 8'h00;
RAM[16'h566B] = 8'h00;
RAM[16'h566C] = 8'h00;
RAM[16'h566D] = 8'h00;
RAM[16'h566E] = 8'h00;
RAM[16'h566F] = 8'h00;
RAM[16'h5670] = 8'h00;
RAM[16'h5671] = 8'h00;
RAM[16'h5672] = 8'h00;
RAM[16'h5673] = 8'h00;
RAM[16'h5674] = 8'h00;
RAM[16'h5675] = 8'h00;
RAM[16'h5676] = 8'h00;
RAM[16'h5677] = 8'h00;
RAM[16'h5678] = 8'h00;
RAM[16'h5679] = 8'h00;
RAM[16'h567A] = 8'h00;
RAM[16'h567B] = 8'h00;
RAM[16'h567C] = 8'h00;
RAM[16'h567D] = 8'h00;
RAM[16'h567E] = 8'h00;
RAM[16'h567F] = 8'h00;
RAM[16'h5680] = 8'h00;
RAM[16'h5681] = 8'h00;
RAM[16'h5682] = 8'h00;
RAM[16'h5683] = 8'h00;
RAM[16'h5684] = 8'h00;
RAM[16'h5685] = 8'h00;
RAM[16'h5686] = 8'h00;
RAM[16'h5687] = 8'h00;
RAM[16'h5688] = 8'h00;
RAM[16'h5689] = 8'h00;
RAM[16'h568A] = 8'h00;
RAM[16'h568B] = 8'h00;
RAM[16'h568C] = 8'h00;
RAM[16'h568D] = 8'h00;
RAM[16'h568E] = 8'h00;
RAM[16'h568F] = 8'h00;
RAM[16'h5690] = 8'h00;
RAM[16'h5691] = 8'h00;
RAM[16'h5692] = 8'h00;
RAM[16'h5693] = 8'h00;
RAM[16'h5694] = 8'h00;
RAM[16'h5695] = 8'h00;
RAM[16'h5696] = 8'h00;
RAM[16'h5697] = 8'h00;
RAM[16'h5698] = 8'h00;
RAM[16'h5699] = 8'h00;
RAM[16'h569A] = 8'h00;
RAM[16'h569B] = 8'h00;
RAM[16'h569C] = 8'h00;
RAM[16'h569D] = 8'h00;
RAM[16'h569E] = 8'h00;
RAM[16'h569F] = 8'h00;
RAM[16'h56A0] = 8'h00;
RAM[16'h56A1] = 8'h00;
RAM[16'h56A2] = 8'h00;
RAM[16'h56A3] = 8'h00;
RAM[16'h56A4] = 8'h00;
RAM[16'h56A5] = 8'h00;
RAM[16'h56A6] = 8'h00;
RAM[16'h56A7] = 8'h00;
RAM[16'h56A8] = 8'h00;
RAM[16'h56A9] = 8'h00;
RAM[16'h56AA] = 8'h00;
RAM[16'h56AB] = 8'h00;
RAM[16'h56AC] = 8'h00;
RAM[16'h56AD] = 8'h00;
RAM[16'h56AE] = 8'h00;
RAM[16'h56AF] = 8'h00;
RAM[16'h56B0] = 8'h00;
RAM[16'h56B1] = 8'h00;
RAM[16'h56B2] = 8'h00;
RAM[16'h56B3] = 8'h00;
RAM[16'h56B4] = 8'h00;
RAM[16'h56B5] = 8'h00;
RAM[16'h56B6] = 8'h00;
RAM[16'h56B7] = 8'h00;
RAM[16'h56B8] = 8'h00;
RAM[16'h56B9] = 8'h00;
RAM[16'h56BA] = 8'h00;
RAM[16'h56BB] = 8'h00;
RAM[16'h56BC] = 8'h00;
RAM[16'h56BD] = 8'h00;
RAM[16'h56BE] = 8'h00;
RAM[16'h56BF] = 8'h00;
RAM[16'h56C0] = 8'h00;
RAM[16'h56C1] = 8'h00;
RAM[16'h56C2] = 8'h00;
RAM[16'h56C3] = 8'h00;
RAM[16'h56C4] = 8'h00;
RAM[16'h56C5] = 8'h00;
RAM[16'h56C6] = 8'h00;
RAM[16'h56C7] = 8'h00;
RAM[16'h56C8] = 8'h00;
RAM[16'h56C9] = 8'h00;
RAM[16'h56CA] = 8'h00;
RAM[16'h56CB] = 8'h00;
RAM[16'h56CC] = 8'h00;
RAM[16'h56CD] = 8'h00;
RAM[16'h56CE] = 8'h00;
RAM[16'h56CF] = 8'h00;
RAM[16'h56D0] = 8'h00;
RAM[16'h56D1] = 8'h00;
RAM[16'h56D2] = 8'h00;
RAM[16'h56D3] = 8'h00;
RAM[16'h56D4] = 8'h00;
RAM[16'h56D5] = 8'h00;
RAM[16'h56D6] = 8'h00;
RAM[16'h56D7] = 8'h00;
RAM[16'h56D8] = 8'h00;
RAM[16'h56D9] = 8'h00;
RAM[16'h56DA] = 8'h00;
RAM[16'h56DB] = 8'h00;
RAM[16'h56DC] = 8'h00;
RAM[16'h56DD] = 8'h00;
RAM[16'h56DE] = 8'h00;
RAM[16'h56DF] = 8'h00;
RAM[16'h56E0] = 8'h00;
RAM[16'h56E1] = 8'h00;
RAM[16'h56E2] = 8'h00;
RAM[16'h56E3] = 8'h00;
RAM[16'h56E4] = 8'h00;
RAM[16'h56E5] = 8'h00;
RAM[16'h56E6] = 8'h00;
RAM[16'h56E7] = 8'h00;
RAM[16'h56E8] = 8'h00;
RAM[16'h56E9] = 8'h00;
RAM[16'h56EA] = 8'h00;
RAM[16'h56EB] = 8'h00;
RAM[16'h56EC] = 8'h00;
RAM[16'h56ED] = 8'h00;
RAM[16'h56EE] = 8'h00;
RAM[16'h56EF] = 8'h00;
RAM[16'h56F0] = 8'h00;
RAM[16'h56F1] = 8'h00;
RAM[16'h56F2] = 8'h00;
RAM[16'h56F3] = 8'h00;
RAM[16'h56F4] = 8'h00;
RAM[16'h56F5] = 8'h00;
RAM[16'h56F6] = 8'h00;
RAM[16'h56F7] = 8'h00;
RAM[16'h56F8] = 8'h00;
RAM[16'h56F9] = 8'h00;
RAM[16'h56FA] = 8'h00;
RAM[16'h56FB] = 8'h00;
RAM[16'h56FC] = 8'h00;
RAM[16'h56FD] = 8'h00;
RAM[16'h56FE] = 8'h00;
RAM[16'h56FF] = 8'h00;
RAM[16'h5700] = 8'h00;
RAM[16'h5701] = 8'h00;
RAM[16'h5702] = 8'h00;
RAM[16'h5703] = 8'h00;
RAM[16'h5704] = 8'h00;
RAM[16'h5705] = 8'h00;
RAM[16'h5706] = 8'h00;
RAM[16'h5707] = 8'h00;
RAM[16'h5708] = 8'h00;
RAM[16'h5709] = 8'h00;
RAM[16'h570A] = 8'h00;
RAM[16'h570B] = 8'h00;
RAM[16'h570C] = 8'h00;
RAM[16'h570D] = 8'h00;
RAM[16'h570E] = 8'h00;
RAM[16'h570F] = 8'h00;
RAM[16'h5710] = 8'h00;
RAM[16'h5711] = 8'h00;
RAM[16'h5712] = 8'h00;
RAM[16'h5713] = 8'h00;
RAM[16'h5714] = 8'h00;
RAM[16'h5715] = 8'h00;
RAM[16'h5716] = 8'h00;
RAM[16'h5717] = 8'h00;
RAM[16'h5718] = 8'h00;
RAM[16'h5719] = 8'h00;
RAM[16'h571A] = 8'h00;
RAM[16'h571B] = 8'h00;
RAM[16'h571C] = 8'h00;
RAM[16'h571D] = 8'h00;
RAM[16'h571E] = 8'h00;
RAM[16'h571F] = 8'h00;
RAM[16'h5720] = 8'h00;
RAM[16'h5721] = 8'h00;
RAM[16'h5722] = 8'h00;
RAM[16'h5723] = 8'h00;
RAM[16'h5724] = 8'h00;
RAM[16'h5725] = 8'h00;
RAM[16'h5726] = 8'h00;
RAM[16'h5727] = 8'h00;
RAM[16'h5728] = 8'h00;
RAM[16'h5729] = 8'h00;
RAM[16'h572A] = 8'h00;
RAM[16'h572B] = 8'h00;
RAM[16'h572C] = 8'h00;
RAM[16'h572D] = 8'h00;
RAM[16'h572E] = 8'h00;
RAM[16'h572F] = 8'h00;
RAM[16'h5730] = 8'h00;
RAM[16'h5731] = 8'h00;
RAM[16'h5732] = 8'h00;
RAM[16'h5733] = 8'h00;
RAM[16'h5734] = 8'h00;
RAM[16'h5735] = 8'h00;
RAM[16'h5736] = 8'h00;
RAM[16'h5737] = 8'h00;
RAM[16'h5738] = 8'h00;
RAM[16'h5739] = 8'h00;
RAM[16'h573A] = 8'h00;
RAM[16'h573B] = 8'h00;
RAM[16'h573C] = 8'h00;
RAM[16'h573D] = 8'h00;
RAM[16'h573E] = 8'h00;
RAM[16'h573F] = 8'h00;
RAM[16'h5740] = 8'h00;
RAM[16'h5741] = 8'h00;
RAM[16'h5742] = 8'h00;
RAM[16'h5743] = 8'h00;
RAM[16'h5744] = 8'h00;
RAM[16'h5745] = 8'h00;
RAM[16'h5746] = 8'h00;
RAM[16'h5747] = 8'h00;
RAM[16'h5748] = 8'h00;
RAM[16'h5749] = 8'h00;
RAM[16'h574A] = 8'h00;
RAM[16'h574B] = 8'h00;
RAM[16'h574C] = 8'h00;
RAM[16'h574D] = 8'h00;
RAM[16'h574E] = 8'h00;
RAM[16'h574F] = 8'h00;
RAM[16'h5750] = 8'h00;
RAM[16'h5751] = 8'h00;
RAM[16'h5752] = 8'h00;
RAM[16'h5753] = 8'h00;
RAM[16'h5754] = 8'h00;
RAM[16'h5755] = 8'h00;
RAM[16'h5756] = 8'h00;
RAM[16'h5757] = 8'h00;
RAM[16'h5758] = 8'h00;
RAM[16'h5759] = 8'h00;
RAM[16'h575A] = 8'h00;
RAM[16'h575B] = 8'h00;
RAM[16'h575C] = 8'h00;
RAM[16'h575D] = 8'h00;
RAM[16'h575E] = 8'h00;
RAM[16'h575F] = 8'h00;
RAM[16'h5760] = 8'h00;
RAM[16'h5761] = 8'h00;
RAM[16'h5762] = 8'h00;
RAM[16'h5763] = 8'h00;
RAM[16'h5764] = 8'h00;
RAM[16'h5765] = 8'h00;
RAM[16'h5766] = 8'h00;
RAM[16'h5767] = 8'h00;
RAM[16'h5768] = 8'h00;
RAM[16'h5769] = 8'h00;
RAM[16'h576A] = 8'h00;
RAM[16'h576B] = 8'h00;
RAM[16'h576C] = 8'h00;
RAM[16'h576D] = 8'h00;
RAM[16'h576E] = 8'h00;
RAM[16'h576F] = 8'h00;
RAM[16'h5770] = 8'h00;
RAM[16'h5771] = 8'h00;
RAM[16'h5772] = 8'h00;
RAM[16'h5773] = 8'h00;
RAM[16'h5774] = 8'h00;
RAM[16'h5775] = 8'h00;
RAM[16'h5776] = 8'h00;
RAM[16'h5777] = 8'h00;
RAM[16'h5778] = 8'h00;
RAM[16'h5779] = 8'h00;
RAM[16'h577A] = 8'h00;
RAM[16'h577B] = 8'h00;
RAM[16'h577C] = 8'h00;
RAM[16'h577D] = 8'h00;
RAM[16'h577E] = 8'h00;
RAM[16'h577F] = 8'h00;
RAM[16'h5780] = 8'h00;
RAM[16'h5781] = 8'h00;
RAM[16'h5782] = 8'h00;
RAM[16'h5783] = 8'h00;
RAM[16'h5784] = 8'h00;
RAM[16'h5785] = 8'h00;
RAM[16'h5786] = 8'h00;
RAM[16'h5787] = 8'h00;
RAM[16'h5788] = 8'h00;
RAM[16'h5789] = 8'h00;
RAM[16'h578A] = 8'h00;
RAM[16'h578B] = 8'h00;
RAM[16'h578C] = 8'h00;
RAM[16'h578D] = 8'h00;
RAM[16'h578E] = 8'h00;
RAM[16'h578F] = 8'h00;
RAM[16'h5790] = 8'h00;
RAM[16'h5791] = 8'h00;
RAM[16'h5792] = 8'h00;
RAM[16'h5793] = 8'h00;
RAM[16'h5794] = 8'h00;
RAM[16'h5795] = 8'h00;
RAM[16'h5796] = 8'h00;
RAM[16'h5797] = 8'h00;
RAM[16'h5798] = 8'h00;
RAM[16'h5799] = 8'h00;
RAM[16'h579A] = 8'h00;
RAM[16'h579B] = 8'h00;
RAM[16'h579C] = 8'h00;
RAM[16'h579D] = 8'h00;
RAM[16'h579E] = 8'h00;
RAM[16'h579F] = 8'h00;
RAM[16'h57A0] = 8'h00;
RAM[16'h57A1] = 8'h00;
RAM[16'h57A2] = 8'h00;
RAM[16'h57A3] = 8'h00;
RAM[16'h57A4] = 8'h00;
RAM[16'h57A5] = 8'h00;
RAM[16'h57A6] = 8'h00;
RAM[16'h57A7] = 8'h00;
RAM[16'h57A8] = 8'h00;
RAM[16'h57A9] = 8'h00;
RAM[16'h57AA] = 8'h00;
RAM[16'h57AB] = 8'h00;
RAM[16'h57AC] = 8'h00;
RAM[16'h57AD] = 8'h00;
RAM[16'h57AE] = 8'h00;
RAM[16'h57AF] = 8'h00;
RAM[16'h57B0] = 8'h00;
RAM[16'h57B1] = 8'h00;
RAM[16'h57B2] = 8'h00;
RAM[16'h57B3] = 8'h00;
RAM[16'h57B4] = 8'h00;
RAM[16'h57B5] = 8'h00;
RAM[16'h57B6] = 8'h00;
RAM[16'h57B7] = 8'h00;
RAM[16'h57B8] = 8'h00;
RAM[16'h57B9] = 8'h00;
RAM[16'h57BA] = 8'h00;
RAM[16'h57BB] = 8'h00;
RAM[16'h57BC] = 8'h00;
RAM[16'h57BD] = 8'h00;
RAM[16'h57BE] = 8'h00;
RAM[16'h57BF] = 8'h00;
RAM[16'h57C0] = 8'h00;
RAM[16'h57C1] = 8'h00;
RAM[16'h57C2] = 8'h00;
RAM[16'h57C3] = 8'h00;
RAM[16'h57C4] = 8'h00;
RAM[16'h57C5] = 8'h00;
RAM[16'h57C6] = 8'h00;
RAM[16'h57C7] = 8'h00;
RAM[16'h57C8] = 8'h00;
RAM[16'h57C9] = 8'h00;
RAM[16'h57CA] = 8'h00;
RAM[16'h57CB] = 8'h00;
RAM[16'h57CC] = 8'h00;
RAM[16'h57CD] = 8'h00;
RAM[16'h57CE] = 8'h00;
RAM[16'h57CF] = 8'h00;
RAM[16'h57D0] = 8'h00;
RAM[16'h57D1] = 8'h00;
RAM[16'h57D2] = 8'h00;
RAM[16'h57D3] = 8'h00;
RAM[16'h57D4] = 8'h00;
RAM[16'h57D5] = 8'h00;
RAM[16'h57D6] = 8'h00;
RAM[16'h57D7] = 8'h00;
RAM[16'h57D8] = 8'h00;
RAM[16'h57D9] = 8'h00;
RAM[16'h57DA] = 8'h00;
RAM[16'h57DB] = 8'h00;
RAM[16'h57DC] = 8'h00;
RAM[16'h57DD] = 8'h00;
RAM[16'h57DE] = 8'h00;
RAM[16'h57DF] = 8'h00;
RAM[16'h57E0] = 8'h00;
RAM[16'h57E1] = 8'h00;
RAM[16'h57E2] = 8'h00;
RAM[16'h57E3] = 8'h00;
RAM[16'h57E4] = 8'h00;
RAM[16'h57E5] = 8'h00;
RAM[16'h57E6] = 8'h00;
RAM[16'h57E7] = 8'h00;
RAM[16'h57E8] = 8'h00;
RAM[16'h57E9] = 8'h00;
RAM[16'h57EA] = 8'h00;
RAM[16'h57EB] = 8'h00;
RAM[16'h57EC] = 8'h00;
RAM[16'h57ED] = 8'h00;
RAM[16'h57EE] = 8'h00;
RAM[16'h57EF] = 8'h00;
RAM[16'h57F0] = 8'h00;
RAM[16'h57F1] = 8'h00;
RAM[16'h57F2] = 8'h00;
RAM[16'h57F3] = 8'h00;
RAM[16'h57F4] = 8'h00;
RAM[16'h57F5] = 8'h00;
RAM[16'h57F6] = 8'h00;
RAM[16'h57F7] = 8'h00;
RAM[16'h57F8] = 8'h00;
RAM[16'h57F9] = 8'h00;
RAM[16'h57FA] = 8'h00;
RAM[16'h57FB] = 8'h00;
RAM[16'h57FC] = 8'h00;
RAM[16'h57FD] = 8'h00;
RAM[16'h57FE] = 8'h00;
RAM[16'h57FF] = 8'h00;
RAM[16'h5800] = 8'h00;
RAM[16'h5801] = 8'h00;
RAM[16'h5802] = 8'h00;
RAM[16'h5803] = 8'h00;
RAM[16'h5804] = 8'h00;
RAM[16'h5805] = 8'h00;
RAM[16'h5806] = 8'h00;
RAM[16'h5807] = 8'h00;
RAM[16'h5808] = 8'h00;
RAM[16'h5809] = 8'h00;
RAM[16'h580A] = 8'h00;
RAM[16'h580B] = 8'h00;
RAM[16'h580C] = 8'h00;
RAM[16'h580D] = 8'h00;
RAM[16'h580E] = 8'h00;
RAM[16'h580F] = 8'h00;
RAM[16'h5810] = 8'h00;
RAM[16'h5811] = 8'h00;
RAM[16'h5812] = 8'h00;
RAM[16'h5813] = 8'h00;
RAM[16'h5814] = 8'h00;
RAM[16'h5815] = 8'h00;
RAM[16'h5816] = 8'h00;
RAM[16'h5817] = 8'h00;
RAM[16'h5818] = 8'h00;
RAM[16'h5819] = 8'h00;
RAM[16'h581A] = 8'h00;
RAM[16'h581B] = 8'h00;
RAM[16'h581C] = 8'h00;
RAM[16'h581D] = 8'h00;
RAM[16'h581E] = 8'h00;
RAM[16'h581F] = 8'h00;
RAM[16'h5820] = 8'h00;
RAM[16'h5821] = 8'h00;
RAM[16'h5822] = 8'h00;
RAM[16'h5823] = 8'h00;
RAM[16'h5824] = 8'h00;
RAM[16'h5825] = 8'h00;
RAM[16'h5826] = 8'h00;
RAM[16'h5827] = 8'h00;
RAM[16'h5828] = 8'h00;
RAM[16'h5829] = 8'h00;
RAM[16'h582A] = 8'h00;
RAM[16'h582B] = 8'h00;
RAM[16'h582C] = 8'h00;
RAM[16'h582D] = 8'h00;
RAM[16'h582E] = 8'h00;
RAM[16'h582F] = 8'h00;
RAM[16'h5830] = 8'h00;
RAM[16'h5831] = 8'h00;
RAM[16'h5832] = 8'h00;
RAM[16'h5833] = 8'h00;
RAM[16'h5834] = 8'h00;
RAM[16'h5835] = 8'h00;
RAM[16'h5836] = 8'h00;
RAM[16'h5837] = 8'h00;
RAM[16'h5838] = 8'h00;
RAM[16'h5839] = 8'h00;
RAM[16'h583A] = 8'h00;
RAM[16'h583B] = 8'h00;
RAM[16'h583C] = 8'h00;
RAM[16'h583D] = 8'h00;
RAM[16'h583E] = 8'h00;
RAM[16'h583F] = 8'h00;
RAM[16'h5840] = 8'h00;
RAM[16'h5841] = 8'h00;
RAM[16'h5842] = 8'h00;
RAM[16'h5843] = 8'h00;
RAM[16'h5844] = 8'h00;
RAM[16'h5845] = 8'h00;
RAM[16'h5846] = 8'h00;
RAM[16'h5847] = 8'h00;
RAM[16'h5848] = 8'h00;
RAM[16'h5849] = 8'h00;
RAM[16'h584A] = 8'h00;
RAM[16'h584B] = 8'h00;
RAM[16'h584C] = 8'h00;
RAM[16'h584D] = 8'h00;
RAM[16'h584E] = 8'h00;
RAM[16'h584F] = 8'h00;
RAM[16'h5850] = 8'h00;
RAM[16'h5851] = 8'h00;
RAM[16'h5852] = 8'h00;
RAM[16'h5853] = 8'h00;
RAM[16'h5854] = 8'h00;
RAM[16'h5855] = 8'h00;
RAM[16'h5856] = 8'h00;
RAM[16'h5857] = 8'h00;
RAM[16'h5858] = 8'h00;
RAM[16'h5859] = 8'h00;
RAM[16'h585A] = 8'h00;
RAM[16'h585B] = 8'h00;
RAM[16'h585C] = 8'h00;
RAM[16'h585D] = 8'h00;
RAM[16'h585E] = 8'h00;
RAM[16'h585F] = 8'h00;
RAM[16'h5860] = 8'h00;
RAM[16'h5861] = 8'h00;
RAM[16'h5862] = 8'h00;
RAM[16'h5863] = 8'h00;
RAM[16'h5864] = 8'h00;
RAM[16'h5865] = 8'h00;
RAM[16'h5866] = 8'h00;
RAM[16'h5867] = 8'h00;
RAM[16'h5868] = 8'h00;
RAM[16'h5869] = 8'h00;
RAM[16'h586A] = 8'h00;
RAM[16'h586B] = 8'h00;
RAM[16'h586C] = 8'h00;
RAM[16'h586D] = 8'h00;
RAM[16'h586E] = 8'h00;
RAM[16'h586F] = 8'h00;
RAM[16'h5870] = 8'h00;
RAM[16'h5871] = 8'h00;
RAM[16'h5872] = 8'h00;
RAM[16'h5873] = 8'h00;
RAM[16'h5874] = 8'h00;
RAM[16'h5875] = 8'h00;
RAM[16'h5876] = 8'h00;
RAM[16'h5877] = 8'h00;
RAM[16'h5878] = 8'h00;
RAM[16'h5879] = 8'h00;
RAM[16'h587A] = 8'h00;
RAM[16'h587B] = 8'h00;
RAM[16'h587C] = 8'h00;
RAM[16'h587D] = 8'h00;
RAM[16'h587E] = 8'h00;
RAM[16'h587F] = 8'h00;
RAM[16'h5880] = 8'h00;
RAM[16'h5881] = 8'h00;
RAM[16'h5882] = 8'h00;
RAM[16'h5883] = 8'h00;
RAM[16'h5884] = 8'h00;
RAM[16'h5885] = 8'h00;
RAM[16'h5886] = 8'h00;
RAM[16'h5887] = 8'h00;
RAM[16'h5888] = 8'h00;
RAM[16'h5889] = 8'h00;
RAM[16'h588A] = 8'h00;
RAM[16'h588B] = 8'h00;
RAM[16'h588C] = 8'h00;
RAM[16'h588D] = 8'h00;
RAM[16'h588E] = 8'h00;
RAM[16'h588F] = 8'h00;
RAM[16'h5890] = 8'h00;
RAM[16'h5891] = 8'h00;
RAM[16'h5892] = 8'h00;
RAM[16'h5893] = 8'h00;
RAM[16'h5894] = 8'h00;
RAM[16'h5895] = 8'h00;
RAM[16'h5896] = 8'h00;
RAM[16'h5897] = 8'h00;
RAM[16'h5898] = 8'h00;
RAM[16'h5899] = 8'h00;
RAM[16'h589A] = 8'h00;
RAM[16'h589B] = 8'h00;
RAM[16'h589C] = 8'h00;
RAM[16'h589D] = 8'h00;
RAM[16'h589E] = 8'h00;
RAM[16'h589F] = 8'h00;
RAM[16'h58A0] = 8'h00;
RAM[16'h58A1] = 8'h00;
RAM[16'h58A2] = 8'h00;
RAM[16'h58A3] = 8'h00;
RAM[16'h58A4] = 8'h00;
RAM[16'h58A5] = 8'h00;
RAM[16'h58A6] = 8'h00;
RAM[16'h58A7] = 8'h00;
RAM[16'h58A8] = 8'h00;
RAM[16'h58A9] = 8'h00;
RAM[16'h58AA] = 8'h00;
RAM[16'h58AB] = 8'h00;
RAM[16'h58AC] = 8'h00;
RAM[16'h58AD] = 8'h00;
RAM[16'h58AE] = 8'h00;
RAM[16'h58AF] = 8'h00;
RAM[16'h58B0] = 8'h00;
RAM[16'h58B1] = 8'h00;
RAM[16'h58B2] = 8'h00;
RAM[16'h58B3] = 8'h00;
RAM[16'h58B4] = 8'h00;
RAM[16'h58B5] = 8'h00;
RAM[16'h58B6] = 8'h00;
RAM[16'h58B7] = 8'h00;
RAM[16'h58B8] = 8'h00;
RAM[16'h58B9] = 8'h00;
RAM[16'h58BA] = 8'h00;
RAM[16'h58BB] = 8'h00;
RAM[16'h58BC] = 8'h00;
RAM[16'h58BD] = 8'h00;
RAM[16'h58BE] = 8'h00;
RAM[16'h58BF] = 8'h00;
RAM[16'h58C0] = 8'h00;
RAM[16'h58C1] = 8'h00;
RAM[16'h58C2] = 8'h00;
RAM[16'h58C3] = 8'h00;
RAM[16'h58C4] = 8'h00;
RAM[16'h58C5] = 8'h00;
RAM[16'h58C6] = 8'h00;
RAM[16'h58C7] = 8'h00;
RAM[16'h58C8] = 8'h00;
RAM[16'h58C9] = 8'h00;
RAM[16'h58CA] = 8'h00;
RAM[16'h58CB] = 8'h00;
RAM[16'h58CC] = 8'h00;
RAM[16'h58CD] = 8'h00;
RAM[16'h58CE] = 8'h00;
RAM[16'h58CF] = 8'h00;
RAM[16'h58D0] = 8'h00;
RAM[16'h58D1] = 8'h00;
RAM[16'h58D2] = 8'h00;
RAM[16'h58D3] = 8'h00;
RAM[16'h58D4] = 8'h00;
RAM[16'h58D5] = 8'h00;
RAM[16'h58D6] = 8'h00;
RAM[16'h58D7] = 8'h00;
RAM[16'h58D8] = 8'h00;
RAM[16'h58D9] = 8'h00;
RAM[16'h58DA] = 8'h00;
RAM[16'h58DB] = 8'h00;
RAM[16'h58DC] = 8'h00;
RAM[16'h58DD] = 8'h00;
RAM[16'h58DE] = 8'h00;
RAM[16'h58DF] = 8'h00;
RAM[16'h58E0] = 8'h00;
RAM[16'h58E1] = 8'h00;
RAM[16'h58E2] = 8'h00;
RAM[16'h58E3] = 8'h00;
RAM[16'h58E4] = 8'h00;
RAM[16'h58E5] = 8'h00;
RAM[16'h58E6] = 8'h00;
RAM[16'h58E7] = 8'h00;
RAM[16'h58E8] = 8'h00;
RAM[16'h58E9] = 8'h00;
RAM[16'h58EA] = 8'h00;
RAM[16'h58EB] = 8'h00;
RAM[16'h58EC] = 8'h00;
RAM[16'h58ED] = 8'h00;
RAM[16'h58EE] = 8'h00;
RAM[16'h58EF] = 8'h00;
RAM[16'h58F0] = 8'h00;
RAM[16'h58F1] = 8'h00;
RAM[16'h58F2] = 8'h00;
RAM[16'h58F3] = 8'h00;
RAM[16'h58F4] = 8'h00;
RAM[16'h58F5] = 8'h00;
RAM[16'h58F6] = 8'h00;
RAM[16'h58F7] = 8'h00;
RAM[16'h58F8] = 8'h00;
RAM[16'h58F9] = 8'h00;
RAM[16'h58FA] = 8'h00;
RAM[16'h58FB] = 8'h00;
RAM[16'h58FC] = 8'h00;
RAM[16'h58FD] = 8'h00;
RAM[16'h58FE] = 8'h00;
RAM[16'h58FF] = 8'h00;
RAM[16'h5900] = 8'h00;
RAM[16'h5901] = 8'h00;
RAM[16'h5902] = 8'h00;
RAM[16'h5903] = 8'h00;
RAM[16'h5904] = 8'h00;
RAM[16'h5905] = 8'h00;
RAM[16'h5906] = 8'h00;
RAM[16'h5907] = 8'h00;
RAM[16'h5908] = 8'h00;
RAM[16'h5909] = 8'h00;
RAM[16'h590A] = 8'h00;
RAM[16'h590B] = 8'h00;
RAM[16'h590C] = 8'h00;
RAM[16'h590D] = 8'h00;
RAM[16'h590E] = 8'h00;
RAM[16'h590F] = 8'h00;
RAM[16'h5910] = 8'h00;
RAM[16'h5911] = 8'h00;
RAM[16'h5912] = 8'h00;
RAM[16'h5913] = 8'h00;
RAM[16'h5914] = 8'h00;
RAM[16'h5915] = 8'h00;
RAM[16'h5916] = 8'h00;
RAM[16'h5917] = 8'h00;
RAM[16'h5918] = 8'h00;
RAM[16'h5919] = 8'h00;
RAM[16'h591A] = 8'h00;
RAM[16'h591B] = 8'h00;
RAM[16'h591C] = 8'h00;
RAM[16'h591D] = 8'h00;
RAM[16'h591E] = 8'h00;
RAM[16'h591F] = 8'h00;
RAM[16'h5920] = 8'h00;
RAM[16'h5921] = 8'h00;
RAM[16'h5922] = 8'h00;
RAM[16'h5923] = 8'h00;
RAM[16'h5924] = 8'h00;
RAM[16'h5925] = 8'h00;
RAM[16'h5926] = 8'h00;
RAM[16'h5927] = 8'h00;
RAM[16'h5928] = 8'h00;
RAM[16'h5929] = 8'h00;
RAM[16'h592A] = 8'h00;
RAM[16'h592B] = 8'h00;
RAM[16'h592C] = 8'h00;
RAM[16'h592D] = 8'h00;
RAM[16'h592E] = 8'h00;
RAM[16'h592F] = 8'h00;
RAM[16'h5930] = 8'h00;
RAM[16'h5931] = 8'h00;
RAM[16'h5932] = 8'h00;
RAM[16'h5933] = 8'h00;
RAM[16'h5934] = 8'h00;
RAM[16'h5935] = 8'h00;
RAM[16'h5936] = 8'h00;
RAM[16'h5937] = 8'h00;
RAM[16'h5938] = 8'h00;
RAM[16'h5939] = 8'h00;
RAM[16'h593A] = 8'h00;
RAM[16'h593B] = 8'h00;
RAM[16'h593C] = 8'h00;
RAM[16'h593D] = 8'h00;
RAM[16'h593E] = 8'h00;
RAM[16'h593F] = 8'h00;
RAM[16'h5940] = 8'h00;
RAM[16'h5941] = 8'h00;
RAM[16'h5942] = 8'h00;
RAM[16'h5943] = 8'h00;
RAM[16'h5944] = 8'h00;
RAM[16'h5945] = 8'h00;
RAM[16'h5946] = 8'h00;
RAM[16'h5947] = 8'h00;
RAM[16'h5948] = 8'h00;
RAM[16'h5949] = 8'h00;
RAM[16'h594A] = 8'h00;
RAM[16'h594B] = 8'h00;
RAM[16'h594C] = 8'h00;
RAM[16'h594D] = 8'h00;
RAM[16'h594E] = 8'h00;
RAM[16'h594F] = 8'h00;
RAM[16'h5950] = 8'h00;
RAM[16'h5951] = 8'h00;
RAM[16'h5952] = 8'h00;
RAM[16'h5953] = 8'h00;
RAM[16'h5954] = 8'h00;
RAM[16'h5955] = 8'h00;
RAM[16'h5956] = 8'h00;
RAM[16'h5957] = 8'h00;
RAM[16'h5958] = 8'h00;
RAM[16'h5959] = 8'h00;
RAM[16'h595A] = 8'h00;
RAM[16'h595B] = 8'h00;
RAM[16'h595C] = 8'h00;
RAM[16'h595D] = 8'h00;
RAM[16'h595E] = 8'h00;
RAM[16'h595F] = 8'h00;
RAM[16'h5960] = 8'h00;
RAM[16'h5961] = 8'h00;
RAM[16'h5962] = 8'h00;
RAM[16'h5963] = 8'h00;
RAM[16'h5964] = 8'h00;
RAM[16'h5965] = 8'h00;
RAM[16'h5966] = 8'h00;
RAM[16'h5967] = 8'h00;
RAM[16'h5968] = 8'h00;
RAM[16'h5969] = 8'h00;
RAM[16'h596A] = 8'h00;
RAM[16'h596B] = 8'h00;
RAM[16'h596C] = 8'h00;
RAM[16'h596D] = 8'h00;
RAM[16'h596E] = 8'h00;
RAM[16'h596F] = 8'h00;
RAM[16'h5970] = 8'h00;
RAM[16'h5971] = 8'h00;
RAM[16'h5972] = 8'h00;
RAM[16'h5973] = 8'h00;
RAM[16'h5974] = 8'h00;
RAM[16'h5975] = 8'h00;
RAM[16'h5976] = 8'h00;
RAM[16'h5977] = 8'h00;
RAM[16'h5978] = 8'h00;
RAM[16'h5979] = 8'h00;
RAM[16'h597A] = 8'h00;
RAM[16'h597B] = 8'h00;
RAM[16'h597C] = 8'h00;
RAM[16'h597D] = 8'h00;
RAM[16'h597E] = 8'h00;
RAM[16'h597F] = 8'h00;
RAM[16'h5980] = 8'h00;
RAM[16'h5981] = 8'h00;
RAM[16'h5982] = 8'h00;
RAM[16'h5983] = 8'h00;
RAM[16'h5984] = 8'h00;
RAM[16'h5985] = 8'h00;
RAM[16'h5986] = 8'h00;
RAM[16'h5987] = 8'h00;
RAM[16'h5988] = 8'h00;
RAM[16'h5989] = 8'h00;
RAM[16'h598A] = 8'h00;
RAM[16'h598B] = 8'h00;
RAM[16'h598C] = 8'h00;
RAM[16'h598D] = 8'h00;
RAM[16'h598E] = 8'h00;
RAM[16'h598F] = 8'h00;
RAM[16'h5990] = 8'h00;
RAM[16'h5991] = 8'h00;
RAM[16'h5992] = 8'h00;
RAM[16'h5993] = 8'h00;
RAM[16'h5994] = 8'h00;
RAM[16'h5995] = 8'h00;
RAM[16'h5996] = 8'h00;
RAM[16'h5997] = 8'h00;
RAM[16'h5998] = 8'h00;
RAM[16'h5999] = 8'h00;
RAM[16'h599A] = 8'h00;
RAM[16'h599B] = 8'h00;
RAM[16'h599C] = 8'h00;
RAM[16'h599D] = 8'h00;
RAM[16'h599E] = 8'h00;
RAM[16'h599F] = 8'h00;
RAM[16'h59A0] = 8'h00;
RAM[16'h59A1] = 8'h00;
RAM[16'h59A2] = 8'h00;
RAM[16'h59A3] = 8'h00;
RAM[16'h59A4] = 8'h00;
RAM[16'h59A5] = 8'h00;
RAM[16'h59A6] = 8'h00;
RAM[16'h59A7] = 8'h00;
RAM[16'h59A8] = 8'h00;
RAM[16'h59A9] = 8'h00;
RAM[16'h59AA] = 8'h00;
RAM[16'h59AB] = 8'h00;
RAM[16'h59AC] = 8'h00;
RAM[16'h59AD] = 8'h00;
RAM[16'h59AE] = 8'h00;
RAM[16'h59AF] = 8'h00;
RAM[16'h59B0] = 8'h00;
RAM[16'h59B1] = 8'h00;
RAM[16'h59B2] = 8'h00;
RAM[16'h59B3] = 8'h00;
RAM[16'h59B4] = 8'h00;
RAM[16'h59B5] = 8'h00;
RAM[16'h59B6] = 8'h00;
RAM[16'h59B7] = 8'h00;
RAM[16'h59B8] = 8'h00;
RAM[16'h59B9] = 8'h00;
RAM[16'h59BA] = 8'h00;
RAM[16'h59BB] = 8'h00;
RAM[16'h59BC] = 8'h00;
RAM[16'h59BD] = 8'h00;
RAM[16'h59BE] = 8'h00;
RAM[16'h59BF] = 8'h00;
RAM[16'h59C0] = 8'h00;
RAM[16'h59C1] = 8'h00;
RAM[16'h59C2] = 8'h00;
RAM[16'h59C3] = 8'h00;
RAM[16'h59C4] = 8'h00;
RAM[16'h59C5] = 8'h00;
RAM[16'h59C6] = 8'h00;
RAM[16'h59C7] = 8'h00;
RAM[16'h59C8] = 8'h00;
RAM[16'h59C9] = 8'h00;
RAM[16'h59CA] = 8'h00;
RAM[16'h59CB] = 8'h00;
RAM[16'h59CC] = 8'h00;
RAM[16'h59CD] = 8'h00;
RAM[16'h59CE] = 8'h00;
RAM[16'h59CF] = 8'h00;
RAM[16'h59D0] = 8'h00;
RAM[16'h59D1] = 8'h00;
RAM[16'h59D2] = 8'h00;
RAM[16'h59D3] = 8'h00;
RAM[16'h59D4] = 8'h00;
RAM[16'h59D5] = 8'h00;
RAM[16'h59D6] = 8'h00;
RAM[16'h59D7] = 8'h00;
RAM[16'h59D8] = 8'h00;
RAM[16'h59D9] = 8'h00;
RAM[16'h59DA] = 8'h00;
RAM[16'h59DB] = 8'h00;
RAM[16'h59DC] = 8'h00;
RAM[16'h59DD] = 8'h00;
RAM[16'h59DE] = 8'h00;
RAM[16'h59DF] = 8'h00;
RAM[16'h59E0] = 8'h00;
RAM[16'h59E1] = 8'h00;
RAM[16'h59E2] = 8'h00;
RAM[16'h59E3] = 8'h00;
RAM[16'h59E4] = 8'h00;
RAM[16'h59E5] = 8'h00;
RAM[16'h59E6] = 8'h00;
RAM[16'h59E7] = 8'h00;
RAM[16'h59E8] = 8'h00;
RAM[16'h59E9] = 8'h00;
RAM[16'h59EA] = 8'h00;
RAM[16'h59EB] = 8'h00;
RAM[16'h59EC] = 8'h00;
RAM[16'h59ED] = 8'h00;
RAM[16'h59EE] = 8'h00;
RAM[16'h59EF] = 8'h00;
RAM[16'h59F0] = 8'h00;
RAM[16'h59F1] = 8'h00;
RAM[16'h59F2] = 8'h00;
RAM[16'h59F3] = 8'h00;
RAM[16'h59F4] = 8'h00;
RAM[16'h59F5] = 8'h00;
RAM[16'h59F6] = 8'h00;
RAM[16'h59F7] = 8'h00;
RAM[16'h59F8] = 8'h00;
RAM[16'h59F9] = 8'h00;
RAM[16'h59FA] = 8'h00;
RAM[16'h59FB] = 8'h00;
RAM[16'h59FC] = 8'h00;
RAM[16'h59FD] = 8'h00;
RAM[16'h59FE] = 8'h00;
RAM[16'h59FF] = 8'h00;
RAM[16'h5A00] = 8'h00;
RAM[16'h5A01] = 8'h00;
RAM[16'h5A02] = 8'h00;
RAM[16'h5A03] = 8'h00;
RAM[16'h5A04] = 8'h00;
RAM[16'h5A05] = 8'h00;
RAM[16'h5A06] = 8'h00;
RAM[16'h5A07] = 8'h00;
RAM[16'h5A08] = 8'h00;
RAM[16'h5A09] = 8'h00;
RAM[16'h5A0A] = 8'h00;
RAM[16'h5A0B] = 8'h00;
RAM[16'h5A0C] = 8'h00;
RAM[16'h5A0D] = 8'h00;
RAM[16'h5A0E] = 8'h00;
RAM[16'h5A0F] = 8'h00;
RAM[16'h5A10] = 8'h00;
RAM[16'h5A11] = 8'h00;
RAM[16'h5A12] = 8'h00;
RAM[16'h5A13] = 8'h00;
RAM[16'h5A14] = 8'h00;
RAM[16'h5A15] = 8'h00;
RAM[16'h5A16] = 8'h00;
RAM[16'h5A17] = 8'h00;
RAM[16'h5A18] = 8'h00;
RAM[16'h5A19] = 8'h00;
RAM[16'h5A1A] = 8'h00;
RAM[16'h5A1B] = 8'h00;
RAM[16'h5A1C] = 8'h00;
RAM[16'h5A1D] = 8'h00;
RAM[16'h5A1E] = 8'h00;
RAM[16'h5A1F] = 8'h00;
RAM[16'h5A20] = 8'h00;
RAM[16'h5A21] = 8'h00;
RAM[16'h5A22] = 8'h00;
RAM[16'h5A23] = 8'h00;
RAM[16'h5A24] = 8'h00;
RAM[16'h5A25] = 8'h00;
RAM[16'h5A26] = 8'h00;
RAM[16'h5A27] = 8'h00;
RAM[16'h5A28] = 8'h00;
RAM[16'h5A29] = 8'h00;
RAM[16'h5A2A] = 8'h00;
RAM[16'h5A2B] = 8'h00;
RAM[16'h5A2C] = 8'h00;
RAM[16'h5A2D] = 8'h00;
RAM[16'h5A2E] = 8'h00;
RAM[16'h5A2F] = 8'h00;
RAM[16'h5A30] = 8'h00;
RAM[16'h5A31] = 8'h00;
RAM[16'h5A32] = 8'h00;
RAM[16'h5A33] = 8'h00;
RAM[16'h5A34] = 8'h00;
RAM[16'h5A35] = 8'h00;
RAM[16'h5A36] = 8'h00;
RAM[16'h5A37] = 8'h00;
RAM[16'h5A38] = 8'h00;
RAM[16'h5A39] = 8'h00;
RAM[16'h5A3A] = 8'h00;
RAM[16'h5A3B] = 8'h00;
RAM[16'h5A3C] = 8'h00;
RAM[16'h5A3D] = 8'h00;
RAM[16'h5A3E] = 8'h00;
RAM[16'h5A3F] = 8'h00;
RAM[16'h5A40] = 8'h00;
RAM[16'h5A41] = 8'h00;
RAM[16'h5A42] = 8'h00;
RAM[16'h5A43] = 8'h00;
RAM[16'h5A44] = 8'h00;
RAM[16'h5A45] = 8'h00;
RAM[16'h5A46] = 8'h00;
RAM[16'h5A47] = 8'h00;
RAM[16'h5A48] = 8'h00;
RAM[16'h5A49] = 8'h00;
RAM[16'h5A4A] = 8'h00;
RAM[16'h5A4B] = 8'h00;
RAM[16'h5A4C] = 8'h00;
RAM[16'h5A4D] = 8'h00;
RAM[16'h5A4E] = 8'h00;
RAM[16'h5A4F] = 8'h00;
RAM[16'h5A50] = 8'h00;
RAM[16'h5A51] = 8'h00;
RAM[16'h5A52] = 8'h00;
RAM[16'h5A53] = 8'h00;
RAM[16'h5A54] = 8'h00;
RAM[16'h5A55] = 8'h00;
RAM[16'h5A56] = 8'h00;
RAM[16'h5A57] = 8'h00;
RAM[16'h5A58] = 8'h00;
RAM[16'h5A59] = 8'h00;
RAM[16'h5A5A] = 8'h00;
RAM[16'h5A5B] = 8'h00;
RAM[16'h5A5C] = 8'h00;
RAM[16'h5A5D] = 8'h00;
RAM[16'h5A5E] = 8'h00;
RAM[16'h5A5F] = 8'h00;
RAM[16'h5A60] = 8'h00;
RAM[16'h5A61] = 8'h00;
RAM[16'h5A62] = 8'h00;
RAM[16'h5A63] = 8'h00;
RAM[16'h5A64] = 8'h00;
RAM[16'h5A65] = 8'h00;
RAM[16'h5A66] = 8'h00;
RAM[16'h5A67] = 8'h00;
RAM[16'h5A68] = 8'h00;
RAM[16'h5A69] = 8'h00;
RAM[16'h5A6A] = 8'h00;
RAM[16'h5A6B] = 8'h00;
RAM[16'h5A6C] = 8'h00;
RAM[16'h5A6D] = 8'h00;
RAM[16'h5A6E] = 8'h00;
RAM[16'h5A6F] = 8'h00;
RAM[16'h5A70] = 8'h00;
RAM[16'h5A71] = 8'h00;
RAM[16'h5A72] = 8'h00;
RAM[16'h5A73] = 8'h00;
RAM[16'h5A74] = 8'h00;
RAM[16'h5A75] = 8'h00;
RAM[16'h5A76] = 8'h00;
RAM[16'h5A77] = 8'h00;
RAM[16'h5A78] = 8'h00;
RAM[16'h5A79] = 8'h00;
RAM[16'h5A7A] = 8'h00;
RAM[16'h5A7B] = 8'h00;
RAM[16'h5A7C] = 8'h00;
RAM[16'h5A7D] = 8'h00;
RAM[16'h5A7E] = 8'h00;
RAM[16'h5A7F] = 8'h00;
RAM[16'h5A80] = 8'h00;
RAM[16'h5A81] = 8'h00;
RAM[16'h5A82] = 8'h00;
RAM[16'h5A83] = 8'h00;
RAM[16'h5A84] = 8'h00;
RAM[16'h5A85] = 8'h00;
RAM[16'h5A86] = 8'h00;
RAM[16'h5A87] = 8'h00;
RAM[16'h5A88] = 8'h00;
RAM[16'h5A89] = 8'h00;
RAM[16'h5A8A] = 8'h00;
RAM[16'h5A8B] = 8'h00;
RAM[16'h5A8C] = 8'h00;
RAM[16'h5A8D] = 8'h00;
RAM[16'h5A8E] = 8'h00;
RAM[16'h5A8F] = 8'h00;
RAM[16'h5A90] = 8'h00;
RAM[16'h5A91] = 8'h00;
RAM[16'h5A92] = 8'h00;
RAM[16'h5A93] = 8'h00;
RAM[16'h5A94] = 8'h00;
RAM[16'h5A95] = 8'h00;
RAM[16'h5A96] = 8'h00;
RAM[16'h5A97] = 8'h00;
RAM[16'h5A98] = 8'h00;
RAM[16'h5A99] = 8'h00;
RAM[16'h5A9A] = 8'h00;
RAM[16'h5A9B] = 8'h00;
RAM[16'h5A9C] = 8'h00;
RAM[16'h5A9D] = 8'h00;
RAM[16'h5A9E] = 8'h00;
RAM[16'h5A9F] = 8'h00;
RAM[16'h5AA0] = 8'h00;
RAM[16'h5AA1] = 8'h00;
RAM[16'h5AA2] = 8'h00;
RAM[16'h5AA3] = 8'h00;
RAM[16'h5AA4] = 8'h00;
RAM[16'h5AA5] = 8'h00;
RAM[16'h5AA6] = 8'h00;
RAM[16'h5AA7] = 8'h00;
RAM[16'h5AA8] = 8'h00;
RAM[16'h5AA9] = 8'h00;
RAM[16'h5AAA] = 8'h00;
RAM[16'h5AAB] = 8'h00;
RAM[16'h5AAC] = 8'h00;
RAM[16'h5AAD] = 8'h00;
RAM[16'h5AAE] = 8'h00;
RAM[16'h5AAF] = 8'h00;
RAM[16'h5AB0] = 8'h00;
RAM[16'h5AB1] = 8'h00;
RAM[16'h5AB2] = 8'h00;
RAM[16'h5AB3] = 8'h00;
RAM[16'h5AB4] = 8'h00;
RAM[16'h5AB5] = 8'h00;
RAM[16'h5AB6] = 8'h00;
RAM[16'h5AB7] = 8'h00;
RAM[16'h5AB8] = 8'h00;
RAM[16'h5AB9] = 8'h00;
RAM[16'h5ABA] = 8'h00;
RAM[16'h5ABB] = 8'h00;
RAM[16'h5ABC] = 8'h00;
RAM[16'h5ABD] = 8'h00;
RAM[16'h5ABE] = 8'h00;
RAM[16'h5ABF] = 8'h00;
RAM[16'h5AC0] = 8'h00;
RAM[16'h5AC1] = 8'h00;
RAM[16'h5AC2] = 8'h00;
RAM[16'h5AC3] = 8'h00;
RAM[16'h5AC4] = 8'h00;
RAM[16'h5AC5] = 8'h00;
RAM[16'h5AC6] = 8'h00;
RAM[16'h5AC7] = 8'h00;
RAM[16'h5AC8] = 8'h00;
RAM[16'h5AC9] = 8'h00;
RAM[16'h5ACA] = 8'h00;
RAM[16'h5ACB] = 8'h00;
RAM[16'h5ACC] = 8'h00;
RAM[16'h5ACD] = 8'h00;
RAM[16'h5ACE] = 8'h00;
RAM[16'h5ACF] = 8'h00;
RAM[16'h5AD0] = 8'h00;
RAM[16'h5AD1] = 8'h00;
RAM[16'h5AD2] = 8'h00;
RAM[16'h5AD3] = 8'h00;
RAM[16'h5AD4] = 8'h00;
RAM[16'h5AD5] = 8'h00;
RAM[16'h5AD6] = 8'h00;
RAM[16'h5AD7] = 8'h00;
RAM[16'h5AD8] = 8'h00;
RAM[16'h5AD9] = 8'h00;
RAM[16'h5ADA] = 8'h00;
RAM[16'h5ADB] = 8'h00;
RAM[16'h5ADC] = 8'h00;
RAM[16'h5ADD] = 8'h00;
RAM[16'h5ADE] = 8'h00;
RAM[16'h5ADF] = 8'h00;
RAM[16'h5AE0] = 8'h00;
RAM[16'h5AE1] = 8'h00;
RAM[16'h5AE2] = 8'h00;
RAM[16'h5AE3] = 8'h00;
RAM[16'h5AE4] = 8'h00;
RAM[16'h5AE5] = 8'h00;
RAM[16'h5AE6] = 8'h00;
RAM[16'h5AE7] = 8'h00;
RAM[16'h5AE8] = 8'h00;
RAM[16'h5AE9] = 8'h00;
RAM[16'h5AEA] = 8'h00;
RAM[16'h5AEB] = 8'h00;
RAM[16'h5AEC] = 8'h00;
RAM[16'h5AED] = 8'h00;
RAM[16'h5AEE] = 8'h00;
RAM[16'h5AEF] = 8'h00;
RAM[16'h5AF0] = 8'h00;
RAM[16'h5AF1] = 8'h00;
RAM[16'h5AF2] = 8'h00;
RAM[16'h5AF3] = 8'h00;
RAM[16'h5AF4] = 8'h00;
RAM[16'h5AF5] = 8'h00;
RAM[16'h5AF6] = 8'h00;
RAM[16'h5AF7] = 8'h00;
RAM[16'h5AF8] = 8'h00;
RAM[16'h5AF9] = 8'h00;
RAM[16'h5AFA] = 8'h00;
RAM[16'h5AFB] = 8'h00;
RAM[16'h5AFC] = 8'h00;
RAM[16'h5AFD] = 8'h00;
RAM[16'h5AFE] = 8'h00;
RAM[16'h5AFF] = 8'h00;
RAM[16'h5B00] = 8'h00;
RAM[16'h5B01] = 8'h00;
RAM[16'h5B02] = 8'h00;
RAM[16'h5B03] = 8'h00;
RAM[16'h5B04] = 8'h00;
RAM[16'h5B05] = 8'h00;
RAM[16'h5B06] = 8'h00;
RAM[16'h5B07] = 8'h00;
RAM[16'h5B08] = 8'h00;
RAM[16'h5B09] = 8'h00;
RAM[16'h5B0A] = 8'h00;
RAM[16'h5B0B] = 8'h00;
RAM[16'h5B0C] = 8'h00;
RAM[16'h5B0D] = 8'h00;
RAM[16'h5B0E] = 8'h00;
RAM[16'h5B0F] = 8'h00;
RAM[16'h5B10] = 8'h00;
RAM[16'h5B11] = 8'h00;
RAM[16'h5B12] = 8'h00;
RAM[16'h5B13] = 8'h00;
RAM[16'h5B14] = 8'h00;
RAM[16'h5B15] = 8'h00;
RAM[16'h5B16] = 8'h00;
RAM[16'h5B17] = 8'h00;
RAM[16'h5B18] = 8'h00;
RAM[16'h5B19] = 8'h00;
RAM[16'h5B1A] = 8'h00;
RAM[16'h5B1B] = 8'h00;
RAM[16'h5B1C] = 8'h00;
RAM[16'h5B1D] = 8'h00;
RAM[16'h5B1E] = 8'h00;
RAM[16'h5B1F] = 8'h00;
RAM[16'h5B20] = 8'h00;
RAM[16'h5B21] = 8'h00;
RAM[16'h5B22] = 8'h00;
RAM[16'h5B23] = 8'h00;
RAM[16'h5B24] = 8'h00;
RAM[16'h5B25] = 8'h00;
RAM[16'h5B26] = 8'h00;
RAM[16'h5B27] = 8'h00;
RAM[16'h5B28] = 8'h00;
RAM[16'h5B29] = 8'h00;
RAM[16'h5B2A] = 8'h00;
RAM[16'h5B2B] = 8'h00;
RAM[16'h5B2C] = 8'h00;
RAM[16'h5B2D] = 8'h00;
RAM[16'h5B2E] = 8'h00;
RAM[16'h5B2F] = 8'h00;
RAM[16'h5B30] = 8'h00;
RAM[16'h5B31] = 8'h00;
RAM[16'h5B32] = 8'h00;
RAM[16'h5B33] = 8'h00;
RAM[16'h5B34] = 8'h00;
RAM[16'h5B35] = 8'h00;
RAM[16'h5B36] = 8'h00;
RAM[16'h5B37] = 8'h00;
RAM[16'h5B38] = 8'h00;
RAM[16'h5B39] = 8'h00;
RAM[16'h5B3A] = 8'h00;
RAM[16'h5B3B] = 8'h00;
RAM[16'h5B3C] = 8'h00;
RAM[16'h5B3D] = 8'h00;
RAM[16'h5B3E] = 8'h00;
RAM[16'h5B3F] = 8'h00;
RAM[16'h5B40] = 8'h00;
RAM[16'h5B41] = 8'h00;
RAM[16'h5B42] = 8'h00;
RAM[16'h5B43] = 8'h00;
RAM[16'h5B44] = 8'h00;
RAM[16'h5B45] = 8'h00;
RAM[16'h5B46] = 8'h00;
RAM[16'h5B47] = 8'h00;
RAM[16'h5B48] = 8'h00;
RAM[16'h5B49] = 8'h00;
RAM[16'h5B4A] = 8'h00;
RAM[16'h5B4B] = 8'h00;
RAM[16'h5B4C] = 8'h00;
RAM[16'h5B4D] = 8'h00;
RAM[16'h5B4E] = 8'h00;
RAM[16'h5B4F] = 8'h00;
RAM[16'h5B50] = 8'h00;
RAM[16'h5B51] = 8'h00;
RAM[16'h5B52] = 8'h00;
RAM[16'h5B53] = 8'h00;
RAM[16'h5B54] = 8'h00;
RAM[16'h5B55] = 8'h00;
RAM[16'h5B56] = 8'h00;
RAM[16'h5B57] = 8'h00;
RAM[16'h5B58] = 8'h00;
RAM[16'h5B59] = 8'h00;
RAM[16'h5B5A] = 8'h00;
RAM[16'h5B5B] = 8'h00;
RAM[16'h5B5C] = 8'h00;
RAM[16'h5B5D] = 8'h00;
RAM[16'h5B5E] = 8'h00;
RAM[16'h5B5F] = 8'h00;
RAM[16'h5B60] = 8'h00;
RAM[16'h5B61] = 8'h00;
RAM[16'h5B62] = 8'h00;
RAM[16'h5B63] = 8'h00;
RAM[16'h5B64] = 8'h00;
RAM[16'h5B65] = 8'h00;
RAM[16'h5B66] = 8'h00;
RAM[16'h5B67] = 8'h00;
RAM[16'h5B68] = 8'h00;
RAM[16'h5B69] = 8'h00;
RAM[16'h5B6A] = 8'h00;
RAM[16'h5B6B] = 8'h00;
RAM[16'h5B6C] = 8'h00;
RAM[16'h5B6D] = 8'h00;
RAM[16'h5B6E] = 8'h00;
RAM[16'h5B6F] = 8'h00;
RAM[16'h5B70] = 8'h00;
RAM[16'h5B71] = 8'h00;
RAM[16'h5B72] = 8'h00;
RAM[16'h5B73] = 8'h00;
RAM[16'h5B74] = 8'h00;
RAM[16'h5B75] = 8'h00;
RAM[16'h5B76] = 8'h00;
RAM[16'h5B77] = 8'h00;
RAM[16'h5B78] = 8'h00;
RAM[16'h5B79] = 8'h00;
RAM[16'h5B7A] = 8'h00;
RAM[16'h5B7B] = 8'h00;
RAM[16'h5B7C] = 8'h00;
RAM[16'h5B7D] = 8'h00;
RAM[16'h5B7E] = 8'h00;
RAM[16'h5B7F] = 8'h00;
RAM[16'h5B80] = 8'h00;
RAM[16'h5B81] = 8'h00;
RAM[16'h5B82] = 8'h00;
RAM[16'h5B83] = 8'h00;
RAM[16'h5B84] = 8'h00;
RAM[16'h5B85] = 8'h00;
RAM[16'h5B86] = 8'h00;
RAM[16'h5B87] = 8'h00;
RAM[16'h5B88] = 8'h00;
RAM[16'h5B89] = 8'h00;
RAM[16'h5B8A] = 8'h00;
RAM[16'h5B8B] = 8'h00;
RAM[16'h5B8C] = 8'h00;
RAM[16'h5B8D] = 8'h00;
RAM[16'h5B8E] = 8'h00;
RAM[16'h5B8F] = 8'h00;
RAM[16'h5B90] = 8'h00;
RAM[16'h5B91] = 8'h00;
RAM[16'h5B92] = 8'h00;
RAM[16'h5B93] = 8'h00;
RAM[16'h5B94] = 8'h00;
RAM[16'h5B95] = 8'h00;
RAM[16'h5B96] = 8'h00;
RAM[16'h5B97] = 8'h00;
RAM[16'h5B98] = 8'h00;
RAM[16'h5B99] = 8'h00;
RAM[16'h5B9A] = 8'h00;
RAM[16'h5B9B] = 8'h00;
RAM[16'h5B9C] = 8'h00;
RAM[16'h5B9D] = 8'h00;
RAM[16'h5B9E] = 8'h00;
RAM[16'h5B9F] = 8'h00;
RAM[16'h5BA0] = 8'h00;
RAM[16'h5BA1] = 8'h00;
RAM[16'h5BA2] = 8'h00;
RAM[16'h5BA3] = 8'h00;
RAM[16'h5BA4] = 8'h00;
RAM[16'h5BA5] = 8'h00;
RAM[16'h5BA6] = 8'h00;
RAM[16'h5BA7] = 8'h00;
RAM[16'h5BA8] = 8'h00;
RAM[16'h5BA9] = 8'h00;
RAM[16'h5BAA] = 8'h00;
RAM[16'h5BAB] = 8'h00;
RAM[16'h5BAC] = 8'h00;
RAM[16'h5BAD] = 8'h00;
RAM[16'h5BAE] = 8'h00;
RAM[16'h5BAF] = 8'h00;
RAM[16'h5BB0] = 8'h00;
RAM[16'h5BB1] = 8'h00;
RAM[16'h5BB2] = 8'h00;
RAM[16'h5BB3] = 8'h00;
RAM[16'h5BB4] = 8'h00;
RAM[16'h5BB5] = 8'h00;
RAM[16'h5BB6] = 8'h00;
RAM[16'h5BB7] = 8'h00;
RAM[16'h5BB8] = 8'h00;
RAM[16'h5BB9] = 8'h00;
RAM[16'h5BBA] = 8'h00;
RAM[16'h5BBB] = 8'h00;
RAM[16'h5BBC] = 8'h00;
RAM[16'h5BBD] = 8'h00;
RAM[16'h5BBE] = 8'h00;
RAM[16'h5BBF] = 8'h00;
RAM[16'h5BC0] = 8'h00;
RAM[16'h5BC1] = 8'h00;
RAM[16'h5BC2] = 8'h00;
RAM[16'h5BC3] = 8'h00;
RAM[16'h5BC4] = 8'h00;
RAM[16'h5BC5] = 8'h00;
RAM[16'h5BC6] = 8'h00;
RAM[16'h5BC7] = 8'h00;
RAM[16'h5BC8] = 8'h00;
RAM[16'h5BC9] = 8'h00;
RAM[16'h5BCA] = 8'h00;
RAM[16'h5BCB] = 8'h00;
RAM[16'h5BCC] = 8'h00;
RAM[16'h5BCD] = 8'h00;
RAM[16'h5BCE] = 8'h00;
RAM[16'h5BCF] = 8'h00;
RAM[16'h5BD0] = 8'h00;
RAM[16'h5BD1] = 8'h00;
RAM[16'h5BD2] = 8'h00;
RAM[16'h5BD3] = 8'h00;
RAM[16'h5BD4] = 8'h00;
RAM[16'h5BD5] = 8'h00;
RAM[16'h5BD6] = 8'h00;
RAM[16'h5BD7] = 8'h00;
RAM[16'h5BD8] = 8'h00;
RAM[16'h5BD9] = 8'h00;
RAM[16'h5BDA] = 8'h00;
RAM[16'h5BDB] = 8'h00;
RAM[16'h5BDC] = 8'h00;
RAM[16'h5BDD] = 8'h00;
RAM[16'h5BDE] = 8'h00;
RAM[16'h5BDF] = 8'h00;
RAM[16'h5BE0] = 8'h00;
RAM[16'h5BE1] = 8'h00;
RAM[16'h5BE2] = 8'h00;
RAM[16'h5BE3] = 8'h00;
RAM[16'h5BE4] = 8'h00;
RAM[16'h5BE5] = 8'h00;
RAM[16'h5BE6] = 8'h00;
RAM[16'h5BE7] = 8'h00;
RAM[16'h5BE8] = 8'h00;
RAM[16'h5BE9] = 8'h00;
RAM[16'h5BEA] = 8'h00;
RAM[16'h5BEB] = 8'h00;
RAM[16'h5BEC] = 8'h00;
RAM[16'h5BED] = 8'h00;
RAM[16'h5BEE] = 8'h00;
RAM[16'h5BEF] = 8'h00;
RAM[16'h5BF0] = 8'h00;
RAM[16'h5BF1] = 8'h00;
RAM[16'h5BF2] = 8'h00;
RAM[16'h5BF3] = 8'h00;
RAM[16'h5BF4] = 8'h00;
RAM[16'h5BF5] = 8'h00;
RAM[16'h5BF6] = 8'h00;
RAM[16'h5BF7] = 8'h00;
RAM[16'h5BF8] = 8'h00;
RAM[16'h5BF9] = 8'h00;
RAM[16'h5BFA] = 8'h00;
RAM[16'h5BFB] = 8'h00;
RAM[16'h5BFC] = 8'h00;
RAM[16'h5BFD] = 8'h00;
RAM[16'h5BFE] = 8'h00;
RAM[16'h5BFF] = 8'h00;
RAM[16'h5C00] = 8'h00;
RAM[16'h5C01] = 8'h00;
RAM[16'h5C02] = 8'h00;
RAM[16'h5C03] = 8'h00;
RAM[16'h5C04] = 8'h00;
RAM[16'h5C05] = 8'h00;
RAM[16'h5C06] = 8'h00;
RAM[16'h5C07] = 8'h00;
RAM[16'h5C08] = 8'h00;
RAM[16'h5C09] = 8'h00;
RAM[16'h5C0A] = 8'h00;
RAM[16'h5C0B] = 8'h00;
RAM[16'h5C0C] = 8'h00;
RAM[16'h5C0D] = 8'h00;
RAM[16'h5C0E] = 8'h00;
RAM[16'h5C0F] = 8'h00;
RAM[16'h5C10] = 8'h00;
RAM[16'h5C11] = 8'h00;
RAM[16'h5C12] = 8'h00;
RAM[16'h5C13] = 8'h00;
RAM[16'h5C14] = 8'h00;
RAM[16'h5C15] = 8'h00;
RAM[16'h5C16] = 8'h00;
RAM[16'h5C17] = 8'h00;
RAM[16'h5C18] = 8'h00;
RAM[16'h5C19] = 8'h00;
RAM[16'h5C1A] = 8'h00;
RAM[16'h5C1B] = 8'h00;
RAM[16'h5C1C] = 8'h00;
RAM[16'h5C1D] = 8'h00;
RAM[16'h5C1E] = 8'h00;
RAM[16'h5C1F] = 8'h00;
RAM[16'h5C20] = 8'h00;
RAM[16'h5C21] = 8'h00;
RAM[16'h5C22] = 8'h00;
RAM[16'h5C23] = 8'h00;
RAM[16'h5C24] = 8'h00;
RAM[16'h5C25] = 8'h00;
RAM[16'h5C26] = 8'h00;
RAM[16'h5C27] = 8'h00;
RAM[16'h5C28] = 8'h00;
RAM[16'h5C29] = 8'h00;
RAM[16'h5C2A] = 8'h00;
RAM[16'h5C2B] = 8'h00;
RAM[16'h5C2C] = 8'h00;
RAM[16'h5C2D] = 8'h00;
RAM[16'h5C2E] = 8'h00;
RAM[16'h5C2F] = 8'h00;
RAM[16'h5C30] = 8'h00;
RAM[16'h5C31] = 8'h00;
RAM[16'h5C32] = 8'h00;
RAM[16'h5C33] = 8'h00;
RAM[16'h5C34] = 8'h00;
RAM[16'h5C35] = 8'h00;
RAM[16'h5C36] = 8'h00;
RAM[16'h5C37] = 8'h00;
RAM[16'h5C38] = 8'h00;
RAM[16'h5C39] = 8'h00;
RAM[16'h5C3A] = 8'h00;
RAM[16'h5C3B] = 8'h00;
RAM[16'h5C3C] = 8'h00;
RAM[16'h5C3D] = 8'h00;
RAM[16'h5C3E] = 8'h00;
RAM[16'h5C3F] = 8'h00;
RAM[16'h5C40] = 8'h00;
RAM[16'h5C41] = 8'h00;
RAM[16'h5C42] = 8'h00;
RAM[16'h5C43] = 8'h00;
RAM[16'h5C44] = 8'h00;
RAM[16'h5C45] = 8'h00;
RAM[16'h5C46] = 8'h00;
RAM[16'h5C47] = 8'h00;
RAM[16'h5C48] = 8'h00;
RAM[16'h5C49] = 8'h00;
RAM[16'h5C4A] = 8'h00;
RAM[16'h5C4B] = 8'h00;
RAM[16'h5C4C] = 8'h00;
RAM[16'h5C4D] = 8'h00;
RAM[16'h5C4E] = 8'h00;
RAM[16'h5C4F] = 8'h00;
RAM[16'h5C50] = 8'h00;
RAM[16'h5C51] = 8'h00;
RAM[16'h5C52] = 8'h00;
RAM[16'h5C53] = 8'h00;
RAM[16'h5C54] = 8'h00;
RAM[16'h5C55] = 8'h00;
RAM[16'h5C56] = 8'h00;
RAM[16'h5C57] = 8'h00;
RAM[16'h5C58] = 8'h00;
RAM[16'h5C59] = 8'h00;
RAM[16'h5C5A] = 8'h00;
RAM[16'h5C5B] = 8'h00;
RAM[16'h5C5C] = 8'h00;
RAM[16'h5C5D] = 8'h00;
RAM[16'h5C5E] = 8'h00;
RAM[16'h5C5F] = 8'h00;
RAM[16'h5C60] = 8'h00;
RAM[16'h5C61] = 8'h00;
RAM[16'h5C62] = 8'h00;
RAM[16'h5C63] = 8'h00;
RAM[16'h5C64] = 8'h00;
RAM[16'h5C65] = 8'h00;
RAM[16'h5C66] = 8'h00;
RAM[16'h5C67] = 8'h00;
RAM[16'h5C68] = 8'h00;
RAM[16'h5C69] = 8'h00;
RAM[16'h5C6A] = 8'h00;
RAM[16'h5C6B] = 8'h00;
RAM[16'h5C6C] = 8'h00;
RAM[16'h5C6D] = 8'h00;
RAM[16'h5C6E] = 8'h00;
RAM[16'h5C6F] = 8'h00;
RAM[16'h5C70] = 8'h00;
RAM[16'h5C71] = 8'h00;
RAM[16'h5C72] = 8'h00;
RAM[16'h5C73] = 8'h00;
RAM[16'h5C74] = 8'h00;
RAM[16'h5C75] = 8'h00;
RAM[16'h5C76] = 8'h00;
RAM[16'h5C77] = 8'h00;
RAM[16'h5C78] = 8'h00;
RAM[16'h5C79] = 8'h00;
RAM[16'h5C7A] = 8'h00;
RAM[16'h5C7B] = 8'h00;
RAM[16'h5C7C] = 8'h00;
RAM[16'h5C7D] = 8'h00;
RAM[16'h5C7E] = 8'h00;
RAM[16'h5C7F] = 8'h00;
RAM[16'h5C80] = 8'h00;
RAM[16'h5C81] = 8'h00;
RAM[16'h5C82] = 8'h00;
RAM[16'h5C83] = 8'h00;
RAM[16'h5C84] = 8'h00;
RAM[16'h5C85] = 8'h00;
RAM[16'h5C86] = 8'h00;
RAM[16'h5C87] = 8'h00;
RAM[16'h5C88] = 8'h00;
RAM[16'h5C89] = 8'h00;
RAM[16'h5C8A] = 8'h00;
RAM[16'h5C8B] = 8'h00;
RAM[16'h5C8C] = 8'h00;
RAM[16'h5C8D] = 8'h00;
RAM[16'h5C8E] = 8'h00;
RAM[16'h5C8F] = 8'h00;
RAM[16'h5C90] = 8'h00;
RAM[16'h5C91] = 8'h00;
RAM[16'h5C92] = 8'h00;
RAM[16'h5C93] = 8'h00;
RAM[16'h5C94] = 8'h00;
RAM[16'h5C95] = 8'h00;
RAM[16'h5C96] = 8'h00;
RAM[16'h5C97] = 8'h00;
RAM[16'h5C98] = 8'h00;
RAM[16'h5C99] = 8'h00;
RAM[16'h5C9A] = 8'h00;
RAM[16'h5C9B] = 8'h00;
RAM[16'h5C9C] = 8'h00;
RAM[16'h5C9D] = 8'h00;
RAM[16'h5C9E] = 8'h00;
RAM[16'h5C9F] = 8'h00;
RAM[16'h5CA0] = 8'h00;
RAM[16'h5CA1] = 8'h00;
RAM[16'h5CA2] = 8'h00;
RAM[16'h5CA3] = 8'h00;
RAM[16'h5CA4] = 8'h00;
RAM[16'h5CA5] = 8'h00;
RAM[16'h5CA6] = 8'h00;
RAM[16'h5CA7] = 8'h00;
RAM[16'h5CA8] = 8'h00;
RAM[16'h5CA9] = 8'h00;
RAM[16'h5CAA] = 8'h00;
RAM[16'h5CAB] = 8'h00;
RAM[16'h5CAC] = 8'h00;
RAM[16'h5CAD] = 8'h00;
RAM[16'h5CAE] = 8'h00;
RAM[16'h5CAF] = 8'h00;
RAM[16'h5CB0] = 8'h00;
RAM[16'h5CB1] = 8'h00;
RAM[16'h5CB2] = 8'h00;
RAM[16'h5CB3] = 8'h00;
RAM[16'h5CB4] = 8'h00;
RAM[16'h5CB5] = 8'h00;
RAM[16'h5CB6] = 8'h00;
RAM[16'h5CB7] = 8'h00;
RAM[16'h5CB8] = 8'h00;
RAM[16'h5CB9] = 8'h00;
RAM[16'h5CBA] = 8'h00;
RAM[16'h5CBB] = 8'h00;
RAM[16'h5CBC] = 8'h00;
RAM[16'h5CBD] = 8'h00;
RAM[16'h5CBE] = 8'h00;
RAM[16'h5CBF] = 8'h00;
RAM[16'h5CC0] = 8'h00;
RAM[16'h5CC1] = 8'h00;
RAM[16'h5CC2] = 8'h00;
RAM[16'h5CC3] = 8'h00;
RAM[16'h5CC4] = 8'h00;
RAM[16'h5CC5] = 8'h00;
RAM[16'h5CC6] = 8'h00;
RAM[16'h5CC7] = 8'h00;
RAM[16'h5CC8] = 8'h00;
RAM[16'h5CC9] = 8'h00;
RAM[16'h5CCA] = 8'h00;
RAM[16'h5CCB] = 8'h00;
RAM[16'h5CCC] = 8'h00;
RAM[16'h5CCD] = 8'h00;
RAM[16'h5CCE] = 8'h00;
RAM[16'h5CCF] = 8'h00;
RAM[16'h5CD0] = 8'h00;
RAM[16'h5CD1] = 8'h00;
RAM[16'h5CD2] = 8'h00;
RAM[16'h5CD3] = 8'h00;
RAM[16'h5CD4] = 8'h00;
RAM[16'h5CD5] = 8'h00;
RAM[16'h5CD6] = 8'h00;
RAM[16'h5CD7] = 8'h00;
RAM[16'h5CD8] = 8'h00;
RAM[16'h5CD9] = 8'h00;
RAM[16'h5CDA] = 8'h00;
RAM[16'h5CDB] = 8'h00;
RAM[16'h5CDC] = 8'h00;
RAM[16'h5CDD] = 8'h00;
RAM[16'h5CDE] = 8'h00;
RAM[16'h5CDF] = 8'h00;
RAM[16'h5CE0] = 8'h00;
RAM[16'h5CE1] = 8'h00;
RAM[16'h5CE2] = 8'h00;
RAM[16'h5CE3] = 8'h00;
RAM[16'h5CE4] = 8'h00;
RAM[16'h5CE5] = 8'h00;
RAM[16'h5CE6] = 8'h00;
RAM[16'h5CE7] = 8'h00;
RAM[16'h5CE8] = 8'h00;
RAM[16'h5CE9] = 8'h00;
RAM[16'h5CEA] = 8'h00;
RAM[16'h5CEB] = 8'h00;
RAM[16'h5CEC] = 8'h00;
RAM[16'h5CED] = 8'h00;
RAM[16'h5CEE] = 8'h00;
RAM[16'h5CEF] = 8'h00;
RAM[16'h5CF0] = 8'h00;
RAM[16'h5CF1] = 8'h00;
RAM[16'h5CF2] = 8'h00;
RAM[16'h5CF3] = 8'h00;
RAM[16'h5CF4] = 8'h00;
RAM[16'h5CF5] = 8'h00;
RAM[16'h5CF6] = 8'h00;
RAM[16'h5CF7] = 8'h00;
RAM[16'h5CF8] = 8'h00;
RAM[16'h5CF9] = 8'h00;
RAM[16'h5CFA] = 8'h00;
RAM[16'h5CFB] = 8'h00;
RAM[16'h5CFC] = 8'h00;
RAM[16'h5CFD] = 8'h00;
RAM[16'h5CFE] = 8'h00;
RAM[16'h5CFF] = 8'h00;
RAM[16'h5D00] = 8'h00;
RAM[16'h5D01] = 8'h00;
RAM[16'h5D02] = 8'h00;
RAM[16'h5D03] = 8'h00;
RAM[16'h5D04] = 8'h00;
RAM[16'h5D05] = 8'h00;
RAM[16'h5D06] = 8'h00;
RAM[16'h5D07] = 8'h00;
RAM[16'h5D08] = 8'h00;
RAM[16'h5D09] = 8'h00;
RAM[16'h5D0A] = 8'h00;
RAM[16'h5D0B] = 8'h00;
RAM[16'h5D0C] = 8'h00;
RAM[16'h5D0D] = 8'h00;
RAM[16'h5D0E] = 8'h00;
RAM[16'h5D0F] = 8'h00;
RAM[16'h5D10] = 8'h00;
RAM[16'h5D11] = 8'h00;
RAM[16'h5D12] = 8'h00;
RAM[16'h5D13] = 8'h00;
RAM[16'h5D14] = 8'h00;
RAM[16'h5D15] = 8'h00;
RAM[16'h5D16] = 8'h00;
RAM[16'h5D17] = 8'h00;
RAM[16'h5D18] = 8'h00;
RAM[16'h5D19] = 8'h00;
RAM[16'h5D1A] = 8'h00;
RAM[16'h5D1B] = 8'h00;
RAM[16'h5D1C] = 8'h00;
RAM[16'h5D1D] = 8'h00;
RAM[16'h5D1E] = 8'h00;
RAM[16'h5D1F] = 8'h00;
RAM[16'h5D20] = 8'h00;
RAM[16'h5D21] = 8'h00;
RAM[16'h5D22] = 8'h00;
RAM[16'h5D23] = 8'h00;
RAM[16'h5D24] = 8'h00;
RAM[16'h5D25] = 8'h00;
RAM[16'h5D26] = 8'h00;
RAM[16'h5D27] = 8'h00;
RAM[16'h5D28] = 8'h00;
RAM[16'h5D29] = 8'h00;
RAM[16'h5D2A] = 8'h00;
RAM[16'h5D2B] = 8'h00;
RAM[16'h5D2C] = 8'h00;
RAM[16'h5D2D] = 8'h00;
RAM[16'h5D2E] = 8'h00;
RAM[16'h5D2F] = 8'h00;
RAM[16'h5D30] = 8'h00;
RAM[16'h5D31] = 8'h00;
RAM[16'h5D32] = 8'h00;
RAM[16'h5D33] = 8'h00;
RAM[16'h5D34] = 8'h00;
RAM[16'h5D35] = 8'h00;
RAM[16'h5D36] = 8'h00;
RAM[16'h5D37] = 8'h00;
RAM[16'h5D38] = 8'h00;
RAM[16'h5D39] = 8'h00;
RAM[16'h5D3A] = 8'h00;
RAM[16'h5D3B] = 8'h00;
RAM[16'h5D3C] = 8'h00;
RAM[16'h5D3D] = 8'h00;
RAM[16'h5D3E] = 8'h00;
RAM[16'h5D3F] = 8'h00;
RAM[16'h5D40] = 8'h00;
RAM[16'h5D41] = 8'h00;
RAM[16'h5D42] = 8'h00;
RAM[16'h5D43] = 8'h00;
RAM[16'h5D44] = 8'h00;
RAM[16'h5D45] = 8'h00;
RAM[16'h5D46] = 8'h00;
RAM[16'h5D47] = 8'h00;
RAM[16'h5D48] = 8'h00;
RAM[16'h5D49] = 8'h00;
RAM[16'h5D4A] = 8'h00;
RAM[16'h5D4B] = 8'h00;
RAM[16'h5D4C] = 8'h00;
RAM[16'h5D4D] = 8'h00;
RAM[16'h5D4E] = 8'h00;
RAM[16'h5D4F] = 8'h00;
RAM[16'h5D50] = 8'h00;
RAM[16'h5D51] = 8'h00;
RAM[16'h5D52] = 8'h00;
RAM[16'h5D53] = 8'h00;
RAM[16'h5D54] = 8'h00;
RAM[16'h5D55] = 8'h00;
RAM[16'h5D56] = 8'h00;
RAM[16'h5D57] = 8'h00;
RAM[16'h5D58] = 8'h00;
RAM[16'h5D59] = 8'h00;
RAM[16'h5D5A] = 8'h00;
RAM[16'h5D5B] = 8'h00;
RAM[16'h5D5C] = 8'h00;
RAM[16'h5D5D] = 8'h00;
RAM[16'h5D5E] = 8'h00;
RAM[16'h5D5F] = 8'h00;
RAM[16'h5D60] = 8'h00;
RAM[16'h5D61] = 8'h00;
RAM[16'h5D62] = 8'h00;
RAM[16'h5D63] = 8'h00;
RAM[16'h5D64] = 8'h00;
RAM[16'h5D65] = 8'h00;
RAM[16'h5D66] = 8'h00;
RAM[16'h5D67] = 8'h00;
RAM[16'h5D68] = 8'h00;
RAM[16'h5D69] = 8'h00;
RAM[16'h5D6A] = 8'h00;
RAM[16'h5D6B] = 8'h00;
RAM[16'h5D6C] = 8'h00;
RAM[16'h5D6D] = 8'h00;
RAM[16'h5D6E] = 8'h00;
RAM[16'h5D6F] = 8'h00;
RAM[16'h5D70] = 8'h00;
RAM[16'h5D71] = 8'h00;
RAM[16'h5D72] = 8'h00;
RAM[16'h5D73] = 8'h00;
RAM[16'h5D74] = 8'h00;
RAM[16'h5D75] = 8'h00;
RAM[16'h5D76] = 8'h00;
RAM[16'h5D77] = 8'h00;
RAM[16'h5D78] = 8'h00;
RAM[16'h5D79] = 8'h00;
RAM[16'h5D7A] = 8'h00;
RAM[16'h5D7B] = 8'h00;
RAM[16'h5D7C] = 8'h00;
RAM[16'h5D7D] = 8'h00;
RAM[16'h5D7E] = 8'h00;
RAM[16'h5D7F] = 8'h00;
RAM[16'h5D80] = 8'h00;
RAM[16'h5D81] = 8'h00;
RAM[16'h5D82] = 8'h00;
RAM[16'h5D83] = 8'h00;
RAM[16'h5D84] = 8'h00;
RAM[16'h5D85] = 8'h00;
RAM[16'h5D86] = 8'h00;
RAM[16'h5D87] = 8'h00;
RAM[16'h5D88] = 8'h00;
RAM[16'h5D89] = 8'h00;
RAM[16'h5D8A] = 8'h00;
RAM[16'h5D8B] = 8'h00;
RAM[16'h5D8C] = 8'h00;
RAM[16'h5D8D] = 8'h00;
RAM[16'h5D8E] = 8'h00;
RAM[16'h5D8F] = 8'h00;
RAM[16'h5D90] = 8'h00;
RAM[16'h5D91] = 8'h00;
RAM[16'h5D92] = 8'h00;
RAM[16'h5D93] = 8'h00;
RAM[16'h5D94] = 8'h00;
RAM[16'h5D95] = 8'h00;
RAM[16'h5D96] = 8'h00;
RAM[16'h5D97] = 8'h00;
RAM[16'h5D98] = 8'h00;
RAM[16'h5D99] = 8'h00;
RAM[16'h5D9A] = 8'h00;
RAM[16'h5D9B] = 8'h00;
RAM[16'h5D9C] = 8'h00;
RAM[16'h5D9D] = 8'h00;
RAM[16'h5D9E] = 8'h00;
RAM[16'h5D9F] = 8'h00;
RAM[16'h5DA0] = 8'h00;
RAM[16'h5DA1] = 8'h00;
RAM[16'h5DA2] = 8'h00;
RAM[16'h5DA3] = 8'h00;
RAM[16'h5DA4] = 8'h00;
RAM[16'h5DA5] = 8'h00;
RAM[16'h5DA6] = 8'h00;
RAM[16'h5DA7] = 8'h00;
RAM[16'h5DA8] = 8'h00;
RAM[16'h5DA9] = 8'h00;
RAM[16'h5DAA] = 8'h00;
RAM[16'h5DAB] = 8'h00;
RAM[16'h5DAC] = 8'h00;
RAM[16'h5DAD] = 8'h00;
RAM[16'h5DAE] = 8'h00;
RAM[16'h5DAF] = 8'h00;
RAM[16'h5DB0] = 8'h00;
RAM[16'h5DB1] = 8'h00;
RAM[16'h5DB2] = 8'h00;
RAM[16'h5DB3] = 8'h00;
RAM[16'h5DB4] = 8'h00;
RAM[16'h5DB5] = 8'h00;
RAM[16'h5DB6] = 8'h00;
RAM[16'h5DB7] = 8'h00;
RAM[16'h5DB8] = 8'h00;
RAM[16'h5DB9] = 8'h00;
RAM[16'h5DBA] = 8'h00;
RAM[16'h5DBB] = 8'h00;
RAM[16'h5DBC] = 8'h00;
RAM[16'h5DBD] = 8'h00;
RAM[16'h5DBE] = 8'h00;
RAM[16'h5DBF] = 8'h00;
RAM[16'h5DC0] = 8'h00;
RAM[16'h5DC1] = 8'h00;
RAM[16'h5DC2] = 8'h00;
RAM[16'h5DC3] = 8'h00;
RAM[16'h5DC4] = 8'h00;
RAM[16'h5DC5] = 8'h00;
RAM[16'h5DC6] = 8'h00;
RAM[16'h5DC7] = 8'h00;
RAM[16'h5DC8] = 8'h00;
RAM[16'h5DC9] = 8'h00;
RAM[16'h5DCA] = 8'h00;
RAM[16'h5DCB] = 8'h00;
RAM[16'h5DCC] = 8'h00;
RAM[16'h5DCD] = 8'h00;
RAM[16'h5DCE] = 8'h00;
RAM[16'h5DCF] = 8'h00;
RAM[16'h5DD0] = 8'h00;
RAM[16'h5DD1] = 8'h00;
RAM[16'h5DD2] = 8'h00;
RAM[16'h5DD3] = 8'h00;
RAM[16'h5DD4] = 8'h00;
RAM[16'h5DD5] = 8'h00;
RAM[16'h5DD6] = 8'h00;
RAM[16'h5DD7] = 8'h00;
RAM[16'h5DD8] = 8'h00;
RAM[16'h5DD9] = 8'h00;
RAM[16'h5DDA] = 8'h00;
RAM[16'h5DDB] = 8'h00;
RAM[16'h5DDC] = 8'h00;
RAM[16'h5DDD] = 8'h00;
RAM[16'h5DDE] = 8'h00;
RAM[16'h5DDF] = 8'h00;
RAM[16'h5DE0] = 8'h00;
RAM[16'h5DE1] = 8'h00;
RAM[16'h5DE2] = 8'h00;
RAM[16'h5DE3] = 8'h00;
RAM[16'h5DE4] = 8'h00;
RAM[16'h5DE5] = 8'h00;
RAM[16'h5DE6] = 8'h00;
RAM[16'h5DE7] = 8'h00;
RAM[16'h5DE8] = 8'h00;
RAM[16'h5DE9] = 8'h00;
RAM[16'h5DEA] = 8'h00;
RAM[16'h5DEB] = 8'h00;
RAM[16'h5DEC] = 8'h00;
RAM[16'h5DED] = 8'h00;
RAM[16'h5DEE] = 8'h00;
RAM[16'h5DEF] = 8'h00;
RAM[16'h5DF0] = 8'h00;
RAM[16'h5DF1] = 8'h00;
RAM[16'h5DF2] = 8'h00;
RAM[16'h5DF3] = 8'h00;
RAM[16'h5DF4] = 8'h00;
RAM[16'h5DF5] = 8'h00;
RAM[16'h5DF6] = 8'h00;
RAM[16'h5DF7] = 8'h00;
RAM[16'h5DF8] = 8'h00;
RAM[16'h5DF9] = 8'h00;
RAM[16'h5DFA] = 8'h00;
RAM[16'h5DFB] = 8'h00;
RAM[16'h5DFC] = 8'h00;
RAM[16'h5DFD] = 8'h00;
RAM[16'h5DFE] = 8'h00;
RAM[16'h5DFF] = 8'h00;
RAM[16'h5E00] = 8'h00;
RAM[16'h5E01] = 8'h00;
RAM[16'h5E02] = 8'h00;
RAM[16'h5E03] = 8'h00;
RAM[16'h5E04] = 8'h00;
RAM[16'h5E05] = 8'h00;
RAM[16'h5E06] = 8'h00;
RAM[16'h5E07] = 8'h00;
RAM[16'h5E08] = 8'h00;
RAM[16'h5E09] = 8'h00;
RAM[16'h5E0A] = 8'h00;
RAM[16'h5E0B] = 8'h00;
RAM[16'h5E0C] = 8'h00;
RAM[16'h5E0D] = 8'h00;
RAM[16'h5E0E] = 8'h00;
RAM[16'h5E0F] = 8'h00;
RAM[16'h5E10] = 8'h00;
RAM[16'h5E11] = 8'h00;
RAM[16'h5E12] = 8'h00;
RAM[16'h5E13] = 8'h00;
RAM[16'h5E14] = 8'h00;
RAM[16'h5E15] = 8'h00;
RAM[16'h5E16] = 8'h00;
RAM[16'h5E17] = 8'h00;
RAM[16'h5E18] = 8'h00;
RAM[16'h5E19] = 8'h00;
RAM[16'h5E1A] = 8'h00;
RAM[16'h5E1B] = 8'h00;
RAM[16'h5E1C] = 8'h00;
RAM[16'h5E1D] = 8'h00;
RAM[16'h5E1E] = 8'h00;
RAM[16'h5E1F] = 8'h00;
RAM[16'h5E20] = 8'h00;
RAM[16'h5E21] = 8'h00;
RAM[16'h5E22] = 8'h00;
RAM[16'h5E23] = 8'h00;
RAM[16'h5E24] = 8'h00;
RAM[16'h5E25] = 8'h00;
RAM[16'h5E26] = 8'h00;
RAM[16'h5E27] = 8'h00;
RAM[16'h5E28] = 8'h00;
RAM[16'h5E29] = 8'h00;
RAM[16'h5E2A] = 8'h00;
RAM[16'h5E2B] = 8'h00;
RAM[16'h5E2C] = 8'h00;
RAM[16'h5E2D] = 8'h00;
RAM[16'h5E2E] = 8'h00;
RAM[16'h5E2F] = 8'h00;
RAM[16'h5E30] = 8'h00;
RAM[16'h5E31] = 8'h00;
RAM[16'h5E32] = 8'h00;
RAM[16'h5E33] = 8'h00;
RAM[16'h5E34] = 8'h00;
RAM[16'h5E35] = 8'h00;
RAM[16'h5E36] = 8'h00;
RAM[16'h5E37] = 8'h00;
RAM[16'h5E38] = 8'h00;
RAM[16'h5E39] = 8'h00;
RAM[16'h5E3A] = 8'h00;
RAM[16'h5E3B] = 8'h00;
RAM[16'h5E3C] = 8'h00;
RAM[16'h5E3D] = 8'h00;
RAM[16'h5E3E] = 8'h00;
RAM[16'h5E3F] = 8'h00;
RAM[16'h5E40] = 8'h00;
RAM[16'h5E41] = 8'h00;
RAM[16'h5E42] = 8'h00;
RAM[16'h5E43] = 8'h00;
RAM[16'h5E44] = 8'h00;
RAM[16'h5E45] = 8'h00;
RAM[16'h5E46] = 8'h00;
RAM[16'h5E47] = 8'h00;
RAM[16'h5E48] = 8'h00;
RAM[16'h5E49] = 8'h00;
RAM[16'h5E4A] = 8'h00;
RAM[16'h5E4B] = 8'h00;
RAM[16'h5E4C] = 8'h00;
RAM[16'h5E4D] = 8'h00;
RAM[16'h5E4E] = 8'h00;
RAM[16'h5E4F] = 8'h00;
RAM[16'h5E50] = 8'h00;
RAM[16'h5E51] = 8'h00;
RAM[16'h5E52] = 8'h00;
RAM[16'h5E53] = 8'h00;
RAM[16'h5E54] = 8'h00;
RAM[16'h5E55] = 8'h00;
RAM[16'h5E56] = 8'h00;
RAM[16'h5E57] = 8'h00;
RAM[16'h5E58] = 8'h00;
RAM[16'h5E59] = 8'h00;
RAM[16'h5E5A] = 8'h00;
RAM[16'h5E5B] = 8'h00;
RAM[16'h5E5C] = 8'h00;
RAM[16'h5E5D] = 8'h00;
RAM[16'h5E5E] = 8'h00;
RAM[16'h5E5F] = 8'h00;
RAM[16'h5E60] = 8'h00;
RAM[16'h5E61] = 8'h00;
RAM[16'h5E62] = 8'h00;
RAM[16'h5E63] = 8'h00;
RAM[16'h5E64] = 8'h00;
RAM[16'h5E65] = 8'h00;
RAM[16'h5E66] = 8'h00;
RAM[16'h5E67] = 8'h00;
RAM[16'h5E68] = 8'h00;
RAM[16'h5E69] = 8'h00;
RAM[16'h5E6A] = 8'h00;
RAM[16'h5E6B] = 8'h00;
RAM[16'h5E6C] = 8'h00;
RAM[16'h5E6D] = 8'h00;
RAM[16'h5E6E] = 8'h00;
RAM[16'h5E6F] = 8'h00;
RAM[16'h5E70] = 8'h00;
RAM[16'h5E71] = 8'h00;
RAM[16'h5E72] = 8'h00;
RAM[16'h5E73] = 8'h00;
RAM[16'h5E74] = 8'h00;
RAM[16'h5E75] = 8'h00;
RAM[16'h5E76] = 8'h00;
RAM[16'h5E77] = 8'h00;
RAM[16'h5E78] = 8'h00;
RAM[16'h5E79] = 8'h00;
RAM[16'h5E7A] = 8'h00;
RAM[16'h5E7B] = 8'h00;
RAM[16'h5E7C] = 8'h00;
RAM[16'h5E7D] = 8'h00;
RAM[16'h5E7E] = 8'h00;
RAM[16'h5E7F] = 8'h00;
RAM[16'h5E80] = 8'h00;
RAM[16'h5E81] = 8'h00;
RAM[16'h5E82] = 8'h00;
RAM[16'h5E83] = 8'h00;
RAM[16'h5E84] = 8'h00;
RAM[16'h5E85] = 8'h00;
RAM[16'h5E86] = 8'h00;
RAM[16'h5E87] = 8'h00;
RAM[16'h5E88] = 8'h00;
RAM[16'h5E89] = 8'h00;
RAM[16'h5E8A] = 8'h00;
RAM[16'h5E8B] = 8'h00;
RAM[16'h5E8C] = 8'h00;
RAM[16'h5E8D] = 8'h00;
RAM[16'h5E8E] = 8'h00;
RAM[16'h5E8F] = 8'h00;
RAM[16'h5E90] = 8'h00;
RAM[16'h5E91] = 8'h00;
RAM[16'h5E92] = 8'h00;
RAM[16'h5E93] = 8'h00;
RAM[16'h5E94] = 8'h00;
RAM[16'h5E95] = 8'h00;
RAM[16'h5E96] = 8'h00;
RAM[16'h5E97] = 8'h00;
RAM[16'h5E98] = 8'h00;
RAM[16'h5E99] = 8'h00;
RAM[16'h5E9A] = 8'h00;
RAM[16'h5E9B] = 8'h00;
RAM[16'h5E9C] = 8'h00;
RAM[16'h5E9D] = 8'h00;
RAM[16'h5E9E] = 8'h00;
RAM[16'h5E9F] = 8'h00;
RAM[16'h5EA0] = 8'h00;
RAM[16'h5EA1] = 8'h00;
RAM[16'h5EA2] = 8'h00;
RAM[16'h5EA3] = 8'h00;
RAM[16'h5EA4] = 8'h00;
RAM[16'h5EA5] = 8'h00;
RAM[16'h5EA6] = 8'h00;
RAM[16'h5EA7] = 8'h00;
RAM[16'h5EA8] = 8'h00;
RAM[16'h5EA9] = 8'h00;
RAM[16'h5EAA] = 8'h00;
RAM[16'h5EAB] = 8'h00;
RAM[16'h5EAC] = 8'h00;
RAM[16'h5EAD] = 8'h00;
RAM[16'h5EAE] = 8'h00;
RAM[16'h5EAF] = 8'h00;
RAM[16'h5EB0] = 8'h00;
RAM[16'h5EB1] = 8'h00;
RAM[16'h5EB2] = 8'h00;
RAM[16'h5EB3] = 8'h00;
RAM[16'h5EB4] = 8'h00;
RAM[16'h5EB5] = 8'h00;
RAM[16'h5EB6] = 8'h00;
RAM[16'h5EB7] = 8'h00;
RAM[16'h5EB8] = 8'h00;
RAM[16'h5EB9] = 8'h00;
RAM[16'h5EBA] = 8'h00;
RAM[16'h5EBB] = 8'h00;
RAM[16'h5EBC] = 8'h00;
RAM[16'h5EBD] = 8'h00;
RAM[16'h5EBE] = 8'h00;
RAM[16'h5EBF] = 8'h00;
RAM[16'h5EC0] = 8'h00;
RAM[16'h5EC1] = 8'h00;
RAM[16'h5EC2] = 8'h00;
RAM[16'h5EC3] = 8'h00;
RAM[16'h5EC4] = 8'h00;
RAM[16'h5EC5] = 8'h00;
RAM[16'h5EC6] = 8'h00;
RAM[16'h5EC7] = 8'h00;
RAM[16'h5EC8] = 8'h00;
RAM[16'h5EC9] = 8'h00;
RAM[16'h5ECA] = 8'h00;
RAM[16'h5ECB] = 8'h00;
RAM[16'h5ECC] = 8'h00;
RAM[16'h5ECD] = 8'h00;
RAM[16'h5ECE] = 8'h00;
RAM[16'h5ECF] = 8'h00;
RAM[16'h5ED0] = 8'h00;
RAM[16'h5ED1] = 8'h00;
RAM[16'h5ED2] = 8'h00;
RAM[16'h5ED3] = 8'h00;
RAM[16'h5ED4] = 8'h00;
RAM[16'h5ED5] = 8'h00;
RAM[16'h5ED6] = 8'h00;
RAM[16'h5ED7] = 8'h00;
RAM[16'h5ED8] = 8'h00;
RAM[16'h5ED9] = 8'h00;
RAM[16'h5EDA] = 8'h00;
RAM[16'h5EDB] = 8'h00;
RAM[16'h5EDC] = 8'h00;
RAM[16'h5EDD] = 8'h00;
RAM[16'h5EDE] = 8'h00;
RAM[16'h5EDF] = 8'h00;
RAM[16'h5EE0] = 8'h00;
RAM[16'h5EE1] = 8'h00;
RAM[16'h5EE2] = 8'h00;
RAM[16'h5EE3] = 8'h00;
RAM[16'h5EE4] = 8'h00;
RAM[16'h5EE5] = 8'h00;
RAM[16'h5EE6] = 8'h00;
RAM[16'h5EE7] = 8'h00;
RAM[16'h5EE8] = 8'h00;
RAM[16'h5EE9] = 8'h00;
RAM[16'h5EEA] = 8'h00;
RAM[16'h5EEB] = 8'h00;
RAM[16'h5EEC] = 8'h00;
RAM[16'h5EED] = 8'h00;
RAM[16'h5EEE] = 8'h00;
RAM[16'h5EEF] = 8'h00;
RAM[16'h5EF0] = 8'h00;
RAM[16'h5EF1] = 8'h00;
RAM[16'h5EF2] = 8'h00;
RAM[16'h5EF3] = 8'h00;
RAM[16'h5EF4] = 8'h00;
RAM[16'h5EF5] = 8'h00;
RAM[16'h5EF6] = 8'h00;
RAM[16'h5EF7] = 8'h00;
RAM[16'h5EF8] = 8'h00;
RAM[16'h5EF9] = 8'h00;
RAM[16'h5EFA] = 8'h00;
RAM[16'h5EFB] = 8'h00;
RAM[16'h5EFC] = 8'h00;
RAM[16'h5EFD] = 8'h00;
RAM[16'h5EFE] = 8'h00;
RAM[16'h5EFF] = 8'h00;
RAM[16'h5F00] = 8'h00;
RAM[16'h5F01] = 8'h00;
RAM[16'h5F02] = 8'h00;
RAM[16'h5F03] = 8'h00;
RAM[16'h5F04] = 8'h00;
RAM[16'h5F05] = 8'h00;
RAM[16'h5F06] = 8'h00;
RAM[16'h5F07] = 8'h00;
RAM[16'h5F08] = 8'h00;
RAM[16'h5F09] = 8'h00;
RAM[16'h5F0A] = 8'h00;
RAM[16'h5F0B] = 8'h00;
RAM[16'h5F0C] = 8'h00;
RAM[16'h5F0D] = 8'h00;
RAM[16'h5F0E] = 8'h00;
RAM[16'h5F0F] = 8'h00;
RAM[16'h5F10] = 8'h00;
RAM[16'h5F11] = 8'h00;
RAM[16'h5F12] = 8'h00;
RAM[16'h5F13] = 8'h00;
RAM[16'h5F14] = 8'h00;
RAM[16'h5F15] = 8'h00;
RAM[16'h5F16] = 8'h00;
RAM[16'h5F17] = 8'h00;
RAM[16'h5F18] = 8'h00;
RAM[16'h5F19] = 8'h00;
RAM[16'h5F1A] = 8'h00;
RAM[16'h5F1B] = 8'h00;
RAM[16'h5F1C] = 8'h00;
RAM[16'h5F1D] = 8'h00;
RAM[16'h5F1E] = 8'h00;
RAM[16'h5F1F] = 8'h00;
RAM[16'h5F20] = 8'h00;
RAM[16'h5F21] = 8'h00;
RAM[16'h5F22] = 8'h00;
RAM[16'h5F23] = 8'h00;
RAM[16'h5F24] = 8'h00;
RAM[16'h5F25] = 8'h00;
RAM[16'h5F26] = 8'h00;
RAM[16'h5F27] = 8'h00;
RAM[16'h5F28] = 8'h00;
RAM[16'h5F29] = 8'h00;
RAM[16'h5F2A] = 8'h00;
RAM[16'h5F2B] = 8'h00;
RAM[16'h5F2C] = 8'h00;
RAM[16'h5F2D] = 8'h00;
RAM[16'h5F2E] = 8'h00;
RAM[16'h5F2F] = 8'h00;
RAM[16'h5F30] = 8'h00;
RAM[16'h5F31] = 8'h00;
RAM[16'h5F32] = 8'h00;
RAM[16'h5F33] = 8'h00;
RAM[16'h5F34] = 8'h00;
RAM[16'h5F35] = 8'h00;
RAM[16'h5F36] = 8'h00;
RAM[16'h5F37] = 8'h00;
RAM[16'h5F38] = 8'h00;
RAM[16'h5F39] = 8'h00;
RAM[16'h5F3A] = 8'h00;
RAM[16'h5F3B] = 8'h00;
RAM[16'h5F3C] = 8'h00;
RAM[16'h5F3D] = 8'h00;
RAM[16'h5F3E] = 8'h00;
RAM[16'h5F3F] = 8'h00;
RAM[16'h5F40] = 8'h00;
RAM[16'h5F41] = 8'h00;
RAM[16'h5F42] = 8'h00;
RAM[16'h5F43] = 8'h00;
RAM[16'h5F44] = 8'h00;
RAM[16'h5F45] = 8'h00;
RAM[16'h5F46] = 8'h00;
RAM[16'h5F47] = 8'h00;
RAM[16'h5F48] = 8'h00;
RAM[16'h5F49] = 8'h00;
RAM[16'h5F4A] = 8'h00;
RAM[16'h5F4B] = 8'h00;
RAM[16'h5F4C] = 8'h00;
RAM[16'h5F4D] = 8'h00;
RAM[16'h5F4E] = 8'h00;
RAM[16'h5F4F] = 8'h00;
RAM[16'h5F50] = 8'h00;
RAM[16'h5F51] = 8'h00;
RAM[16'h5F52] = 8'h00;
RAM[16'h5F53] = 8'h00;
RAM[16'h5F54] = 8'h00;
RAM[16'h5F55] = 8'h00;
RAM[16'h5F56] = 8'h00;
RAM[16'h5F57] = 8'h00;
RAM[16'h5F58] = 8'h00;
RAM[16'h5F59] = 8'h00;
RAM[16'h5F5A] = 8'h00;
RAM[16'h5F5B] = 8'h00;
RAM[16'h5F5C] = 8'h00;
RAM[16'h5F5D] = 8'h00;
RAM[16'h5F5E] = 8'h00;
RAM[16'h5F5F] = 8'h00;
RAM[16'h5F60] = 8'h00;
RAM[16'h5F61] = 8'h00;
RAM[16'h5F62] = 8'h00;
RAM[16'h5F63] = 8'h00;
RAM[16'h5F64] = 8'h00;
RAM[16'h5F65] = 8'h00;
RAM[16'h5F66] = 8'h00;
RAM[16'h5F67] = 8'h00;
RAM[16'h5F68] = 8'h00;
RAM[16'h5F69] = 8'h00;
RAM[16'h5F6A] = 8'h00;
RAM[16'h5F6B] = 8'h00;
RAM[16'h5F6C] = 8'h00;
RAM[16'h5F6D] = 8'h00;
RAM[16'h5F6E] = 8'h00;
RAM[16'h5F6F] = 8'h00;
RAM[16'h5F70] = 8'h00;
RAM[16'h5F71] = 8'h00;
RAM[16'h5F72] = 8'h00;
RAM[16'h5F73] = 8'h00;
RAM[16'h5F74] = 8'h00;
RAM[16'h5F75] = 8'h00;
RAM[16'h5F76] = 8'h00;
RAM[16'h5F77] = 8'h00;
RAM[16'h5F78] = 8'h00;
RAM[16'h5F79] = 8'h00;
RAM[16'h5F7A] = 8'h00;
RAM[16'h5F7B] = 8'h00;
RAM[16'h5F7C] = 8'h00;
RAM[16'h5F7D] = 8'h00;
RAM[16'h5F7E] = 8'h00;
RAM[16'h5F7F] = 8'h00;
RAM[16'h5F80] = 8'h00;
RAM[16'h5F81] = 8'h00;
RAM[16'h5F82] = 8'h00;
RAM[16'h5F83] = 8'h00;
RAM[16'h5F84] = 8'h00;
RAM[16'h5F85] = 8'h00;
RAM[16'h5F86] = 8'h00;
RAM[16'h5F87] = 8'h00;
RAM[16'h5F88] = 8'h00;
RAM[16'h5F89] = 8'h00;
RAM[16'h5F8A] = 8'h00;
RAM[16'h5F8B] = 8'h00;
RAM[16'h5F8C] = 8'h00;
RAM[16'h5F8D] = 8'h00;
RAM[16'h5F8E] = 8'h00;
RAM[16'h5F8F] = 8'h00;
RAM[16'h5F90] = 8'h00;
RAM[16'h5F91] = 8'h00;
RAM[16'h5F92] = 8'h00;
RAM[16'h5F93] = 8'h00;
RAM[16'h5F94] = 8'h00;
RAM[16'h5F95] = 8'h00;
RAM[16'h5F96] = 8'h00;
RAM[16'h5F97] = 8'h00;
RAM[16'h5F98] = 8'h00;
RAM[16'h5F99] = 8'h00;
RAM[16'h5F9A] = 8'h00;
RAM[16'h5F9B] = 8'h00;
RAM[16'h5F9C] = 8'h00;
RAM[16'h5F9D] = 8'h00;
RAM[16'h5F9E] = 8'h00;
RAM[16'h5F9F] = 8'h00;
RAM[16'h5FA0] = 8'h00;
RAM[16'h5FA1] = 8'h00;
RAM[16'h5FA2] = 8'h00;
RAM[16'h5FA3] = 8'h00;
RAM[16'h5FA4] = 8'h00;
RAM[16'h5FA5] = 8'h00;
RAM[16'h5FA6] = 8'h00;
RAM[16'h5FA7] = 8'h00;
RAM[16'h5FA8] = 8'h00;
RAM[16'h5FA9] = 8'h00;
RAM[16'h5FAA] = 8'h00;
RAM[16'h5FAB] = 8'h00;
RAM[16'h5FAC] = 8'h00;
RAM[16'h5FAD] = 8'h00;
RAM[16'h5FAE] = 8'h00;
RAM[16'h5FAF] = 8'h00;
RAM[16'h5FB0] = 8'h00;
RAM[16'h5FB1] = 8'h00;
RAM[16'h5FB2] = 8'h00;
RAM[16'h5FB3] = 8'h00;
RAM[16'h5FB4] = 8'h00;
RAM[16'h5FB5] = 8'h00;
RAM[16'h5FB6] = 8'h00;
RAM[16'h5FB7] = 8'h00;
RAM[16'h5FB8] = 8'h00;
RAM[16'h5FB9] = 8'h00;
RAM[16'h5FBA] = 8'h00;
RAM[16'h5FBB] = 8'h00;
RAM[16'h5FBC] = 8'h00;
RAM[16'h5FBD] = 8'h00;
RAM[16'h5FBE] = 8'h00;
RAM[16'h5FBF] = 8'h00;
RAM[16'h5FC0] = 8'h00;
RAM[16'h5FC1] = 8'h00;
RAM[16'h5FC2] = 8'h00;
RAM[16'h5FC3] = 8'h00;
RAM[16'h5FC4] = 8'h00;
RAM[16'h5FC5] = 8'h00;
RAM[16'h5FC6] = 8'h00;
RAM[16'h5FC7] = 8'h00;
RAM[16'h5FC8] = 8'h00;
RAM[16'h5FC9] = 8'h00;
RAM[16'h5FCA] = 8'h00;
RAM[16'h5FCB] = 8'h00;
RAM[16'h5FCC] = 8'h00;
RAM[16'h5FCD] = 8'h00;
RAM[16'h5FCE] = 8'h00;
RAM[16'h5FCF] = 8'h00;
RAM[16'h5FD0] = 8'h00;
RAM[16'h5FD1] = 8'h00;
RAM[16'h5FD2] = 8'h00;
RAM[16'h5FD3] = 8'h00;
RAM[16'h5FD4] = 8'h00;
RAM[16'h5FD5] = 8'h00;
RAM[16'h5FD6] = 8'h00;
RAM[16'h5FD7] = 8'h00;
RAM[16'h5FD8] = 8'h00;
RAM[16'h5FD9] = 8'h00;
RAM[16'h5FDA] = 8'h00;
RAM[16'h5FDB] = 8'h00;
RAM[16'h5FDC] = 8'h00;
RAM[16'h5FDD] = 8'h00;
RAM[16'h5FDE] = 8'h00;
RAM[16'h5FDF] = 8'h00;
RAM[16'h5FE0] = 8'h00;
RAM[16'h5FE1] = 8'h00;
RAM[16'h5FE2] = 8'h00;
RAM[16'h5FE3] = 8'h00;
RAM[16'h5FE4] = 8'h00;
RAM[16'h5FE5] = 8'h00;
RAM[16'h5FE6] = 8'h00;
RAM[16'h5FE7] = 8'h00;
RAM[16'h5FE8] = 8'h00;
RAM[16'h5FE9] = 8'h00;
RAM[16'h5FEA] = 8'h00;
RAM[16'h5FEB] = 8'h00;
RAM[16'h5FEC] = 8'h00;
RAM[16'h5FED] = 8'h00;
RAM[16'h5FEE] = 8'h00;
RAM[16'h5FEF] = 8'h00;
RAM[16'h5FF0] = 8'h00;
RAM[16'h5FF1] = 8'h00;
RAM[16'h5FF2] = 8'h00;
RAM[16'h5FF3] = 8'h00;
RAM[16'h5FF4] = 8'h00;
RAM[16'h5FF5] = 8'h00;
RAM[16'h5FF6] = 8'h00;
RAM[16'h5FF7] = 8'h00;
RAM[16'h5FF8] = 8'h00;
RAM[16'h5FF9] = 8'h00;
RAM[16'h5FFA] = 8'h00;
RAM[16'h5FFB] = 8'h00;
RAM[16'h5FFC] = 8'h00;
RAM[16'h5FFD] = 8'h00;
RAM[16'h5FFE] = 8'h00;
RAM[16'h5FFF] = 8'h00;
RAM[16'h6000] = 8'h00;
RAM[16'h6001] = 8'h00;
RAM[16'h6002] = 8'h00;
RAM[16'h6003] = 8'h00;
RAM[16'h6004] = 8'h00;
RAM[16'h6005] = 8'h00;
RAM[16'h6006] = 8'h00;
RAM[16'h6007] = 8'h00;
RAM[16'h6008] = 8'h00;
RAM[16'h6009] = 8'h00;
RAM[16'h600A] = 8'h00;
RAM[16'h600B] = 8'h00;
RAM[16'h600C] = 8'h00;
RAM[16'h600D] = 8'h00;
RAM[16'h600E] = 8'h00;
RAM[16'h600F] = 8'h00;
RAM[16'h6010] = 8'h00;
RAM[16'h6011] = 8'h00;
RAM[16'h6012] = 8'h00;
RAM[16'h6013] = 8'h00;
RAM[16'h6014] = 8'h00;
RAM[16'h6015] = 8'h00;
RAM[16'h6016] = 8'h00;
RAM[16'h6017] = 8'h00;
RAM[16'h6018] = 8'h00;
RAM[16'h6019] = 8'h00;
RAM[16'h601A] = 8'h00;
RAM[16'h601B] = 8'h00;
RAM[16'h601C] = 8'h00;
RAM[16'h601D] = 8'h00;
RAM[16'h601E] = 8'h00;
RAM[16'h601F] = 8'h00;
RAM[16'h6020] = 8'h00;
RAM[16'h6021] = 8'h00;
RAM[16'h6022] = 8'h00;
RAM[16'h6023] = 8'h00;
RAM[16'h6024] = 8'h00;
RAM[16'h6025] = 8'h00;
RAM[16'h6026] = 8'h00;
RAM[16'h6027] = 8'h00;
RAM[16'h6028] = 8'h00;
RAM[16'h6029] = 8'h00;
RAM[16'h602A] = 8'h00;
RAM[16'h602B] = 8'h00;
RAM[16'h602C] = 8'h00;
RAM[16'h602D] = 8'h00;
RAM[16'h602E] = 8'h00;
RAM[16'h602F] = 8'h00;
RAM[16'h6030] = 8'h00;
RAM[16'h6031] = 8'h00;
RAM[16'h6032] = 8'h00;
RAM[16'h6033] = 8'h00;
RAM[16'h6034] = 8'h00;
RAM[16'h6035] = 8'h00;
RAM[16'h6036] = 8'h00;
RAM[16'h6037] = 8'h00;
RAM[16'h6038] = 8'h00;
RAM[16'h6039] = 8'h00;
RAM[16'h603A] = 8'h00;
RAM[16'h603B] = 8'h00;
RAM[16'h603C] = 8'h00;
RAM[16'h603D] = 8'h00;
RAM[16'h603E] = 8'h00;
RAM[16'h603F] = 8'h00;
RAM[16'h6040] = 8'h00;
RAM[16'h6041] = 8'h00;
RAM[16'h6042] = 8'h00;
RAM[16'h6043] = 8'h00;
RAM[16'h6044] = 8'h00;
RAM[16'h6045] = 8'h00;
RAM[16'h6046] = 8'h00;
RAM[16'h6047] = 8'h00;
RAM[16'h6048] = 8'h00;
RAM[16'h6049] = 8'h00;
RAM[16'h604A] = 8'h00;
RAM[16'h604B] = 8'h00;
RAM[16'h604C] = 8'h00;
RAM[16'h604D] = 8'h00;
RAM[16'h604E] = 8'h00;
RAM[16'h604F] = 8'h00;
RAM[16'h6050] = 8'h00;
RAM[16'h6051] = 8'h00;
RAM[16'h6052] = 8'h00;
RAM[16'h6053] = 8'h00;
RAM[16'h6054] = 8'h00;
RAM[16'h6055] = 8'h00;
RAM[16'h6056] = 8'h00;
RAM[16'h6057] = 8'h00;
RAM[16'h6058] = 8'h00;
RAM[16'h6059] = 8'h00;
RAM[16'h605A] = 8'h00;
RAM[16'h605B] = 8'h00;
RAM[16'h605C] = 8'h00;
RAM[16'h605D] = 8'h00;
RAM[16'h605E] = 8'h00;
RAM[16'h605F] = 8'h00;
RAM[16'h6060] = 8'h00;
RAM[16'h6061] = 8'h00;
RAM[16'h6062] = 8'h00;
RAM[16'h6063] = 8'h00;
RAM[16'h6064] = 8'h00;
RAM[16'h6065] = 8'h00;
RAM[16'h6066] = 8'h00;
RAM[16'h6067] = 8'h00;
RAM[16'h6068] = 8'h00;
RAM[16'h6069] = 8'h00;
RAM[16'h606A] = 8'h00;
RAM[16'h606B] = 8'h00;
RAM[16'h606C] = 8'h00;
RAM[16'h606D] = 8'h00;
RAM[16'h606E] = 8'h00;
RAM[16'h606F] = 8'h00;
RAM[16'h6070] = 8'h00;
RAM[16'h6071] = 8'h00;
RAM[16'h6072] = 8'h00;
RAM[16'h6073] = 8'h00;
RAM[16'h6074] = 8'h00;
RAM[16'h6075] = 8'h00;
RAM[16'h6076] = 8'h00;
RAM[16'h6077] = 8'h00;
RAM[16'h6078] = 8'h00;
RAM[16'h6079] = 8'h00;
RAM[16'h607A] = 8'h00;
RAM[16'h607B] = 8'h00;
RAM[16'h607C] = 8'h00;
RAM[16'h607D] = 8'h00;
RAM[16'h607E] = 8'h00;
RAM[16'h607F] = 8'h00;
RAM[16'h6080] = 8'h00;
RAM[16'h6081] = 8'h00;
RAM[16'h6082] = 8'h00;
RAM[16'h6083] = 8'h00;
RAM[16'h6084] = 8'h00;
RAM[16'h6085] = 8'h00;
RAM[16'h6086] = 8'h00;
RAM[16'h6087] = 8'h00;
RAM[16'h6088] = 8'h00;
RAM[16'h6089] = 8'h00;
RAM[16'h608A] = 8'h00;
RAM[16'h608B] = 8'h00;
RAM[16'h608C] = 8'h00;
RAM[16'h608D] = 8'h00;
RAM[16'h608E] = 8'h00;
RAM[16'h608F] = 8'h00;
RAM[16'h6090] = 8'h00;
RAM[16'h6091] = 8'h00;
RAM[16'h6092] = 8'h00;
RAM[16'h6093] = 8'h00;
RAM[16'h6094] = 8'h00;
RAM[16'h6095] = 8'h00;
RAM[16'h6096] = 8'h00;
RAM[16'h6097] = 8'h00;
RAM[16'h6098] = 8'h00;
RAM[16'h6099] = 8'h00;
RAM[16'h609A] = 8'h00;
RAM[16'h609B] = 8'h00;
RAM[16'h609C] = 8'h00;
RAM[16'h609D] = 8'h00;
RAM[16'h609E] = 8'h00;
RAM[16'h609F] = 8'h00;
RAM[16'h60A0] = 8'h00;
RAM[16'h60A1] = 8'h00;
RAM[16'h60A2] = 8'h00;
RAM[16'h60A3] = 8'h00;
RAM[16'h60A4] = 8'h00;
RAM[16'h60A5] = 8'h00;
RAM[16'h60A6] = 8'h00;
RAM[16'h60A7] = 8'h00;
RAM[16'h60A8] = 8'h00;
RAM[16'h60A9] = 8'h00;
RAM[16'h60AA] = 8'h00;
RAM[16'h60AB] = 8'h00;
RAM[16'h60AC] = 8'h00;
RAM[16'h60AD] = 8'h00;
RAM[16'h60AE] = 8'h00;
RAM[16'h60AF] = 8'h00;
RAM[16'h60B0] = 8'h00;
RAM[16'h60B1] = 8'h00;
RAM[16'h60B2] = 8'h00;
RAM[16'h60B3] = 8'h00;
RAM[16'h60B4] = 8'h00;
RAM[16'h60B5] = 8'h00;
RAM[16'h60B6] = 8'h00;
RAM[16'h60B7] = 8'h00;
RAM[16'h60B8] = 8'h00;
RAM[16'h60B9] = 8'h00;
RAM[16'h60BA] = 8'h00;
RAM[16'h60BB] = 8'h00;
RAM[16'h60BC] = 8'h00;
RAM[16'h60BD] = 8'h00;
RAM[16'h60BE] = 8'h00;
RAM[16'h60BF] = 8'h00;
RAM[16'h60C0] = 8'h00;
RAM[16'h60C1] = 8'h00;
RAM[16'h60C2] = 8'h00;
RAM[16'h60C3] = 8'h00;
RAM[16'h60C4] = 8'h00;
RAM[16'h60C5] = 8'h00;
RAM[16'h60C6] = 8'h00;
RAM[16'h60C7] = 8'h00;
RAM[16'h60C8] = 8'h00;
RAM[16'h60C9] = 8'h00;
RAM[16'h60CA] = 8'h00;
RAM[16'h60CB] = 8'h00;
RAM[16'h60CC] = 8'h00;
RAM[16'h60CD] = 8'h00;
RAM[16'h60CE] = 8'h00;
RAM[16'h60CF] = 8'h00;
RAM[16'h60D0] = 8'h00;
RAM[16'h60D1] = 8'h00;
RAM[16'h60D2] = 8'h00;
RAM[16'h60D3] = 8'h00;
RAM[16'h60D4] = 8'h00;
RAM[16'h60D5] = 8'h00;
RAM[16'h60D6] = 8'h00;
RAM[16'h60D7] = 8'h00;
RAM[16'h60D8] = 8'h00;
RAM[16'h60D9] = 8'h00;
RAM[16'h60DA] = 8'h00;
RAM[16'h60DB] = 8'h00;
RAM[16'h60DC] = 8'h00;
RAM[16'h60DD] = 8'h00;
RAM[16'h60DE] = 8'h00;
RAM[16'h60DF] = 8'h00;
RAM[16'h60E0] = 8'h00;
RAM[16'h60E1] = 8'h00;
RAM[16'h60E2] = 8'h00;
RAM[16'h60E3] = 8'h00;
RAM[16'h60E4] = 8'h00;
RAM[16'h60E5] = 8'h00;
RAM[16'h60E6] = 8'h00;
RAM[16'h60E7] = 8'h00;
RAM[16'h60E8] = 8'h00;
RAM[16'h60E9] = 8'h00;
RAM[16'h60EA] = 8'h00;
RAM[16'h60EB] = 8'h00;
RAM[16'h60EC] = 8'h00;
RAM[16'h60ED] = 8'h00;
RAM[16'h60EE] = 8'h00;
RAM[16'h60EF] = 8'h00;
RAM[16'h60F0] = 8'h00;
RAM[16'h60F1] = 8'h00;
RAM[16'h60F2] = 8'h00;
RAM[16'h60F3] = 8'h00;
RAM[16'h60F4] = 8'h00;
RAM[16'h60F5] = 8'h00;
RAM[16'h60F6] = 8'h00;
RAM[16'h60F7] = 8'h00;
RAM[16'h60F8] = 8'h00;
RAM[16'h60F9] = 8'h00;
RAM[16'h60FA] = 8'h00;
RAM[16'h60FB] = 8'h00;
RAM[16'h60FC] = 8'h00;
RAM[16'h60FD] = 8'h00;
RAM[16'h60FE] = 8'h00;
RAM[16'h60FF] = 8'h00;
RAM[16'h6100] = 8'h00;
RAM[16'h6101] = 8'h00;
RAM[16'h6102] = 8'h00;
RAM[16'h6103] = 8'h00;
RAM[16'h6104] = 8'h00;
RAM[16'h6105] = 8'h00;
RAM[16'h6106] = 8'h00;
RAM[16'h6107] = 8'h00;
RAM[16'h6108] = 8'h00;
RAM[16'h6109] = 8'h00;
RAM[16'h610A] = 8'h00;
RAM[16'h610B] = 8'h00;
RAM[16'h610C] = 8'h00;
RAM[16'h610D] = 8'h00;
RAM[16'h610E] = 8'h00;
RAM[16'h610F] = 8'h00;
RAM[16'h6110] = 8'h00;
RAM[16'h6111] = 8'h00;
RAM[16'h6112] = 8'h00;
RAM[16'h6113] = 8'h00;
RAM[16'h6114] = 8'h00;
RAM[16'h6115] = 8'h00;
RAM[16'h6116] = 8'h00;
RAM[16'h6117] = 8'h00;
RAM[16'h6118] = 8'h00;
RAM[16'h6119] = 8'h00;
RAM[16'h611A] = 8'h00;
RAM[16'h611B] = 8'h00;
RAM[16'h611C] = 8'h00;
RAM[16'h611D] = 8'h00;
RAM[16'h611E] = 8'h00;
RAM[16'h611F] = 8'h00;
RAM[16'h6120] = 8'h00;
RAM[16'h6121] = 8'h00;
RAM[16'h6122] = 8'h00;
RAM[16'h6123] = 8'h00;
RAM[16'h6124] = 8'h00;
RAM[16'h6125] = 8'h00;
RAM[16'h6126] = 8'h00;
RAM[16'h6127] = 8'h00;
RAM[16'h6128] = 8'h00;
RAM[16'h6129] = 8'h00;
RAM[16'h612A] = 8'h00;
RAM[16'h612B] = 8'h00;
RAM[16'h612C] = 8'h00;
RAM[16'h612D] = 8'h00;
RAM[16'h612E] = 8'h00;
RAM[16'h612F] = 8'h00;
RAM[16'h6130] = 8'h00;
RAM[16'h6131] = 8'h00;
RAM[16'h6132] = 8'h00;
RAM[16'h6133] = 8'h00;
RAM[16'h6134] = 8'h00;
RAM[16'h6135] = 8'h00;
RAM[16'h6136] = 8'h00;
RAM[16'h6137] = 8'h00;
RAM[16'h6138] = 8'h00;
RAM[16'h6139] = 8'h00;
RAM[16'h613A] = 8'h00;
RAM[16'h613B] = 8'h00;
RAM[16'h613C] = 8'h00;
RAM[16'h613D] = 8'h00;
RAM[16'h613E] = 8'h00;
RAM[16'h613F] = 8'h00;
RAM[16'h6140] = 8'h00;
RAM[16'h6141] = 8'h00;
RAM[16'h6142] = 8'h00;
RAM[16'h6143] = 8'h00;
RAM[16'h6144] = 8'h00;
RAM[16'h6145] = 8'h00;
RAM[16'h6146] = 8'h00;
RAM[16'h6147] = 8'h00;
RAM[16'h6148] = 8'h00;
RAM[16'h6149] = 8'h00;
RAM[16'h614A] = 8'h00;
RAM[16'h614B] = 8'h00;
RAM[16'h614C] = 8'h00;
RAM[16'h614D] = 8'h00;
RAM[16'h614E] = 8'h00;
RAM[16'h614F] = 8'h00;
RAM[16'h6150] = 8'h00;
RAM[16'h6151] = 8'h00;
RAM[16'h6152] = 8'h00;
RAM[16'h6153] = 8'h00;
RAM[16'h6154] = 8'h00;
RAM[16'h6155] = 8'h00;
RAM[16'h6156] = 8'h00;
RAM[16'h6157] = 8'h00;
RAM[16'h6158] = 8'h00;
RAM[16'h6159] = 8'h00;
RAM[16'h615A] = 8'h00;
RAM[16'h615B] = 8'h00;
RAM[16'h615C] = 8'h00;
RAM[16'h615D] = 8'h00;
RAM[16'h615E] = 8'h00;
RAM[16'h615F] = 8'h00;
RAM[16'h6160] = 8'h00;
RAM[16'h6161] = 8'h00;
RAM[16'h6162] = 8'h00;
RAM[16'h6163] = 8'h00;
RAM[16'h6164] = 8'h00;
RAM[16'h6165] = 8'h00;
RAM[16'h6166] = 8'h00;
RAM[16'h6167] = 8'h00;
RAM[16'h6168] = 8'h00;
RAM[16'h6169] = 8'h00;
RAM[16'h616A] = 8'h00;
RAM[16'h616B] = 8'h00;
RAM[16'h616C] = 8'h00;
RAM[16'h616D] = 8'h00;
RAM[16'h616E] = 8'h00;
RAM[16'h616F] = 8'h00;
RAM[16'h6170] = 8'h00;
RAM[16'h6171] = 8'h00;
RAM[16'h6172] = 8'h00;
RAM[16'h6173] = 8'h00;
RAM[16'h6174] = 8'h00;
RAM[16'h6175] = 8'h00;
RAM[16'h6176] = 8'h00;
RAM[16'h6177] = 8'h00;
RAM[16'h6178] = 8'h00;
RAM[16'h6179] = 8'h00;
RAM[16'h617A] = 8'h00;
RAM[16'h617B] = 8'h00;
RAM[16'h617C] = 8'h00;
RAM[16'h617D] = 8'h00;
RAM[16'h617E] = 8'h00;
RAM[16'h617F] = 8'h00;
RAM[16'h6180] = 8'h00;
RAM[16'h6181] = 8'h00;
RAM[16'h6182] = 8'h00;
RAM[16'h6183] = 8'h00;
RAM[16'h6184] = 8'h00;
RAM[16'h6185] = 8'h00;
RAM[16'h6186] = 8'h00;
RAM[16'h6187] = 8'h00;
RAM[16'h6188] = 8'h00;
RAM[16'h6189] = 8'h00;
RAM[16'h618A] = 8'h00;
RAM[16'h618B] = 8'h00;
RAM[16'h618C] = 8'h00;
RAM[16'h618D] = 8'h00;
RAM[16'h618E] = 8'h00;
RAM[16'h618F] = 8'h00;
RAM[16'h6190] = 8'h00;
RAM[16'h6191] = 8'h00;
RAM[16'h6192] = 8'h00;
RAM[16'h6193] = 8'h00;
RAM[16'h6194] = 8'h00;
RAM[16'h6195] = 8'h00;
RAM[16'h6196] = 8'h00;
RAM[16'h6197] = 8'h00;
RAM[16'h6198] = 8'h00;
RAM[16'h6199] = 8'h00;
RAM[16'h619A] = 8'h00;
RAM[16'h619B] = 8'h00;
RAM[16'h619C] = 8'h00;
RAM[16'h619D] = 8'h00;
RAM[16'h619E] = 8'h00;
RAM[16'h619F] = 8'h00;
RAM[16'h61A0] = 8'h00;
RAM[16'h61A1] = 8'h00;
RAM[16'h61A2] = 8'h00;
RAM[16'h61A3] = 8'h00;
RAM[16'h61A4] = 8'h00;
RAM[16'h61A5] = 8'h00;
RAM[16'h61A6] = 8'h00;
RAM[16'h61A7] = 8'h00;
RAM[16'h61A8] = 8'h00;
RAM[16'h61A9] = 8'h00;
RAM[16'h61AA] = 8'h00;
RAM[16'h61AB] = 8'h00;
RAM[16'h61AC] = 8'h00;
RAM[16'h61AD] = 8'h00;
RAM[16'h61AE] = 8'h00;
RAM[16'h61AF] = 8'h00;
RAM[16'h61B0] = 8'h00;
RAM[16'h61B1] = 8'h00;
RAM[16'h61B2] = 8'h00;
RAM[16'h61B3] = 8'h00;
RAM[16'h61B4] = 8'h00;
RAM[16'h61B5] = 8'h00;
RAM[16'h61B6] = 8'h00;
RAM[16'h61B7] = 8'h00;
RAM[16'h61B8] = 8'h00;
RAM[16'h61B9] = 8'h00;
RAM[16'h61BA] = 8'h00;
RAM[16'h61BB] = 8'h00;
RAM[16'h61BC] = 8'h00;
RAM[16'h61BD] = 8'h00;
RAM[16'h61BE] = 8'h00;
RAM[16'h61BF] = 8'h00;
RAM[16'h61C0] = 8'h00;
RAM[16'h61C1] = 8'h00;
RAM[16'h61C2] = 8'h00;
RAM[16'h61C3] = 8'h00;
RAM[16'h61C4] = 8'h00;
RAM[16'h61C5] = 8'h00;
RAM[16'h61C6] = 8'h00;
RAM[16'h61C7] = 8'h00;
RAM[16'h61C8] = 8'h00;
RAM[16'h61C9] = 8'h00;
RAM[16'h61CA] = 8'h00;
RAM[16'h61CB] = 8'h00;
RAM[16'h61CC] = 8'h00;
RAM[16'h61CD] = 8'h00;
RAM[16'h61CE] = 8'h00;
RAM[16'h61CF] = 8'h00;
RAM[16'h61D0] = 8'h00;
RAM[16'h61D1] = 8'h00;
RAM[16'h61D2] = 8'h00;
RAM[16'h61D3] = 8'h00;
RAM[16'h61D4] = 8'h00;
RAM[16'h61D5] = 8'h00;
RAM[16'h61D6] = 8'h00;
RAM[16'h61D7] = 8'h00;
RAM[16'h61D8] = 8'h00;
RAM[16'h61D9] = 8'h00;
RAM[16'h61DA] = 8'h00;
RAM[16'h61DB] = 8'h00;
RAM[16'h61DC] = 8'h00;
RAM[16'h61DD] = 8'h00;
RAM[16'h61DE] = 8'h00;
RAM[16'h61DF] = 8'h00;
RAM[16'h61E0] = 8'h00;
RAM[16'h61E1] = 8'h00;
RAM[16'h61E2] = 8'h00;
RAM[16'h61E3] = 8'h00;
RAM[16'h61E4] = 8'h00;
RAM[16'h61E5] = 8'h00;
RAM[16'h61E6] = 8'h00;
RAM[16'h61E7] = 8'h00;
RAM[16'h61E8] = 8'h00;
RAM[16'h61E9] = 8'h00;
RAM[16'h61EA] = 8'h00;
RAM[16'h61EB] = 8'h00;
RAM[16'h61EC] = 8'h00;
RAM[16'h61ED] = 8'h00;
RAM[16'h61EE] = 8'h00;
RAM[16'h61EF] = 8'h00;
RAM[16'h61F0] = 8'h00;
RAM[16'h61F1] = 8'h00;
RAM[16'h61F2] = 8'h00;
RAM[16'h61F3] = 8'h00;
RAM[16'h61F4] = 8'h00;
RAM[16'h61F5] = 8'h00;
RAM[16'h61F6] = 8'h00;
RAM[16'h61F7] = 8'h00;
RAM[16'h61F8] = 8'h00;
RAM[16'h61F9] = 8'h00;
RAM[16'h61FA] = 8'h00;
RAM[16'h61FB] = 8'h00;
RAM[16'h61FC] = 8'h00;
RAM[16'h61FD] = 8'h00;
RAM[16'h61FE] = 8'h00;
RAM[16'h61FF] = 8'h00;
RAM[16'h6200] = 8'h00;
RAM[16'h6201] = 8'h00;
RAM[16'h6202] = 8'h00;
RAM[16'h6203] = 8'h00;
RAM[16'h6204] = 8'h00;
RAM[16'h6205] = 8'h00;
RAM[16'h6206] = 8'h00;
RAM[16'h6207] = 8'h00;
RAM[16'h6208] = 8'h00;
RAM[16'h6209] = 8'h00;
RAM[16'h620A] = 8'h00;
RAM[16'h620B] = 8'h00;
RAM[16'h620C] = 8'h00;
RAM[16'h620D] = 8'h00;
RAM[16'h620E] = 8'h00;
RAM[16'h620F] = 8'h00;
RAM[16'h6210] = 8'h00;
RAM[16'h6211] = 8'h00;
RAM[16'h6212] = 8'h00;
RAM[16'h6213] = 8'h00;
RAM[16'h6214] = 8'h00;
RAM[16'h6215] = 8'h00;
RAM[16'h6216] = 8'h00;
RAM[16'h6217] = 8'h00;
RAM[16'h6218] = 8'h00;
RAM[16'h6219] = 8'h00;
RAM[16'h621A] = 8'h00;
RAM[16'h621B] = 8'h00;
RAM[16'h621C] = 8'h00;
RAM[16'h621D] = 8'h00;
RAM[16'h621E] = 8'h00;
RAM[16'h621F] = 8'h00;
RAM[16'h6220] = 8'h00;
RAM[16'h6221] = 8'h00;
RAM[16'h6222] = 8'h00;
RAM[16'h6223] = 8'h00;
RAM[16'h6224] = 8'h00;
RAM[16'h6225] = 8'h00;
RAM[16'h6226] = 8'h00;
RAM[16'h6227] = 8'h00;
RAM[16'h6228] = 8'h00;
RAM[16'h6229] = 8'h00;
RAM[16'h622A] = 8'h00;
RAM[16'h622B] = 8'h00;
RAM[16'h622C] = 8'h00;
RAM[16'h622D] = 8'h00;
RAM[16'h622E] = 8'h00;
RAM[16'h622F] = 8'h00;
RAM[16'h6230] = 8'h00;
RAM[16'h6231] = 8'h00;
RAM[16'h6232] = 8'h00;
RAM[16'h6233] = 8'h00;
RAM[16'h6234] = 8'h00;
RAM[16'h6235] = 8'h00;
RAM[16'h6236] = 8'h00;
RAM[16'h6237] = 8'h00;
RAM[16'h6238] = 8'h00;
RAM[16'h6239] = 8'h00;
RAM[16'h623A] = 8'h00;
RAM[16'h623B] = 8'h00;
RAM[16'h623C] = 8'h00;
RAM[16'h623D] = 8'h00;
RAM[16'h623E] = 8'h00;
RAM[16'h623F] = 8'h00;
RAM[16'h6240] = 8'h00;
RAM[16'h6241] = 8'h00;
RAM[16'h6242] = 8'h00;
RAM[16'h6243] = 8'h00;
RAM[16'h6244] = 8'h00;
RAM[16'h6245] = 8'h00;
RAM[16'h6246] = 8'h00;
RAM[16'h6247] = 8'h00;
RAM[16'h6248] = 8'h00;
RAM[16'h6249] = 8'h00;
RAM[16'h624A] = 8'h00;
RAM[16'h624B] = 8'h00;
RAM[16'h624C] = 8'h00;
RAM[16'h624D] = 8'h00;
RAM[16'h624E] = 8'h00;
RAM[16'h624F] = 8'h00;
RAM[16'h6250] = 8'h00;
RAM[16'h6251] = 8'h00;
RAM[16'h6252] = 8'h00;
RAM[16'h6253] = 8'h00;
RAM[16'h6254] = 8'h00;
RAM[16'h6255] = 8'h00;
RAM[16'h6256] = 8'h00;
RAM[16'h6257] = 8'h00;
RAM[16'h6258] = 8'h00;
RAM[16'h6259] = 8'h00;
RAM[16'h625A] = 8'h00;
RAM[16'h625B] = 8'h00;
RAM[16'h625C] = 8'h00;
RAM[16'h625D] = 8'h00;
RAM[16'h625E] = 8'h00;
RAM[16'h625F] = 8'h00;
RAM[16'h6260] = 8'h00;
RAM[16'h6261] = 8'h00;
RAM[16'h6262] = 8'h00;
RAM[16'h6263] = 8'h00;
RAM[16'h6264] = 8'h00;
RAM[16'h6265] = 8'h00;
RAM[16'h6266] = 8'h00;
RAM[16'h6267] = 8'h00;
RAM[16'h6268] = 8'h00;
RAM[16'h6269] = 8'h00;
RAM[16'h626A] = 8'h00;
RAM[16'h626B] = 8'h00;
RAM[16'h626C] = 8'h00;
RAM[16'h626D] = 8'h00;
RAM[16'h626E] = 8'h00;
RAM[16'h626F] = 8'h00;
RAM[16'h6270] = 8'h00;
RAM[16'h6271] = 8'h00;
RAM[16'h6272] = 8'h00;
RAM[16'h6273] = 8'h00;
RAM[16'h6274] = 8'h00;
RAM[16'h6275] = 8'h00;
RAM[16'h6276] = 8'h00;
RAM[16'h6277] = 8'h00;
RAM[16'h6278] = 8'h00;
RAM[16'h6279] = 8'h00;
RAM[16'h627A] = 8'h00;
RAM[16'h627B] = 8'h00;
RAM[16'h627C] = 8'h00;
RAM[16'h627D] = 8'h00;
RAM[16'h627E] = 8'h00;
RAM[16'h627F] = 8'h00;
RAM[16'h6280] = 8'h00;
RAM[16'h6281] = 8'h00;
RAM[16'h6282] = 8'h00;
RAM[16'h6283] = 8'h00;
RAM[16'h6284] = 8'h00;
RAM[16'h6285] = 8'h00;
RAM[16'h6286] = 8'h00;
RAM[16'h6287] = 8'h00;
RAM[16'h6288] = 8'h00;
RAM[16'h6289] = 8'h00;
RAM[16'h628A] = 8'h00;
RAM[16'h628B] = 8'h00;
RAM[16'h628C] = 8'h00;
RAM[16'h628D] = 8'h00;
RAM[16'h628E] = 8'h00;
RAM[16'h628F] = 8'h00;
RAM[16'h6290] = 8'h00;
RAM[16'h6291] = 8'h00;
RAM[16'h6292] = 8'h00;
RAM[16'h6293] = 8'h00;
RAM[16'h6294] = 8'h00;
RAM[16'h6295] = 8'h00;
RAM[16'h6296] = 8'h00;
RAM[16'h6297] = 8'h00;
RAM[16'h6298] = 8'h00;
RAM[16'h6299] = 8'h00;
RAM[16'h629A] = 8'h00;
RAM[16'h629B] = 8'h00;
RAM[16'h629C] = 8'h00;
RAM[16'h629D] = 8'h00;
RAM[16'h629E] = 8'h00;
RAM[16'h629F] = 8'h00;
RAM[16'h62A0] = 8'h00;
RAM[16'h62A1] = 8'h00;
RAM[16'h62A2] = 8'h00;
RAM[16'h62A3] = 8'h00;
RAM[16'h62A4] = 8'h00;
RAM[16'h62A5] = 8'h00;
RAM[16'h62A6] = 8'h00;
RAM[16'h62A7] = 8'h00;
RAM[16'h62A8] = 8'h00;
RAM[16'h62A9] = 8'h00;
RAM[16'h62AA] = 8'h00;
RAM[16'h62AB] = 8'h00;
RAM[16'h62AC] = 8'h00;
RAM[16'h62AD] = 8'h00;
RAM[16'h62AE] = 8'h00;
RAM[16'h62AF] = 8'h00;
RAM[16'h62B0] = 8'h00;
RAM[16'h62B1] = 8'h00;
RAM[16'h62B2] = 8'h00;
RAM[16'h62B3] = 8'h00;
RAM[16'h62B4] = 8'h00;
RAM[16'h62B5] = 8'h00;
RAM[16'h62B6] = 8'h00;
RAM[16'h62B7] = 8'h00;
RAM[16'h62B8] = 8'h00;
RAM[16'h62B9] = 8'h00;
RAM[16'h62BA] = 8'h00;
RAM[16'h62BB] = 8'h00;
RAM[16'h62BC] = 8'h00;
RAM[16'h62BD] = 8'h00;
RAM[16'h62BE] = 8'h00;
RAM[16'h62BF] = 8'h00;
RAM[16'h62C0] = 8'h00;
RAM[16'h62C1] = 8'h00;
RAM[16'h62C2] = 8'h00;
RAM[16'h62C3] = 8'h00;
RAM[16'h62C4] = 8'h00;
RAM[16'h62C5] = 8'h00;
RAM[16'h62C6] = 8'h00;
RAM[16'h62C7] = 8'h00;
RAM[16'h62C8] = 8'h00;
RAM[16'h62C9] = 8'h00;
RAM[16'h62CA] = 8'h00;
RAM[16'h62CB] = 8'h00;
RAM[16'h62CC] = 8'h00;
RAM[16'h62CD] = 8'h00;
RAM[16'h62CE] = 8'h00;
RAM[16'h62CF] = 8'h00;
RAM[16'h62D0] = 8'h00;
RAM[16'h62D1] = 8'h00;
RAM[16'h62D2] = 8'h00;
RAM[16'h62D3] = 8'h00;
RAM[16'h62D4] = 8'h00;
RAM[16'h62D5] = 8'h00;
RAM[16'h62D6] = 8'h00;
RAM[16'h62D7] = 8'h00;
RAM[16'h62D8] = 8'h00;
RAM[16'h62D9] = 8'h00;
RAM[16'h62DA] = 8'h00;
RAM[16'h62DB] = 8'h00;
RAM[16'h62DC] = 8'h00;
RAM[16'h62DD] = 8'h00;
RAM[16'h62DE] = 8'h00;
RAM[16'h62DF] = 8'h00;
RAM[16'h62E0] = 8'h00;
RAM[16'h62E1] = 8'h00;
RAM[16'h62E2] = 8'h00;
RAM[16'h62E3] = 8'h00;
RAM[16'h62E4] = 8'h00;
RAM[16'h62E5] = 8'h00;
RAM[16'h62E6] = 8'h00;
RAM[16'h62E7] = 8'h00;
RAM[16'h62E8] = 8'h00;
RAM[16'h62E9] = 8'h00;
RAM[16'h62EA] = 8'h00;
RAM[16'h62EB] = 8'h00;
RAM[16'h62EC] = 8'h00;
RAM[16'h62ED] = 8'h00;
RAM[16'h62EE] = 8'h00;
RAM[16'h62EF] = 8'h00;
RAM[16'h62F0] = 8'h00;
RAM[16'h62F1] = 8'h00;
RAM[16'h62F2] = 8'h00;
RAM[16'h62F3] = 8'h00;
RAM[16'h62F4] = 8'h00;
RAM[16'h62F5] = 8'h00;
RAM[16'h62F6] = 8'h00;
RAM[16'h62F7] = 8'h00;
RAM[16'h62F8] = 8'h00;
RAM[16'h62F9] = 8'h00;
RAM[16'h62FA] = 8'h00;
RAM[16'h62FB] = 8'h00;
RAM[16'h62FC] = 8'h00;
RAM[16'h62FD] = 8'h00;
RAM[16'h62FE] = 8'h00;
RAM[16'h62FF] = 8'h00;
RAM[16'h6300] = 8'h00;
RAM[16'h6301] = 8'h00;
RAM[16'h6302] = 8'h00;
RAM[16'h6303] = 8'h00;
RAM[16'h6304] = 8'h00;
RAM[16'h6305] = 8'h00;
RAM[16'h6306] = 8'h00;
RAM[16'h6307] = 8'h00;
RAM[16'h6308] = 8'h00;
RAM[16'h6309] = 8'h00;
RAM[16'h630A] = 8'h00;
RAM[16'h630B] = 8'h00;
RAM[16'h630C] = 8'h00;
RAM[16'h630D] = 8'h00;
RAM[16'h630E] = 8'h00;
RAM[16'h630F] = 8'h00;
RAM[16'h6310] = 8'h00;
RAM[16'h6311] = 8'h00;
RAM[16'h6312] = 8'h00;
RAM[16'h6313] = 8'h00;
RAM[16'h6314] = 8'h00;
RAM[16'h6315] = 8'h00;
RAM[16'h6316] = 8'h00;
RAM[16'h6317] = 8'h00;
RAM[16'h6318] = 8'h00;
RAM[16'h6319] = 8'h00;
RAM[16'h631A] = 8'h00;
RAM[16'h631B] = 8'h00;
RAM[16'h631C] = 8'h00;
RAM[16'h631D] = 8'h00;
RAM[16'h631E] = 8'h00;
RAM[16'h631F] = 8'h00;
RAM[16'h6320] = 8'h00;
RAM[16'h6321] = 8'h00;
RAM[16'h6322] = 8'h00;
RAM[16'h6323] = 8'h00;
RAM[16'h6324] = 8'h00;
RAM[16'h6325] = 8'h00;
RAM[16'h6326] = 8'h00;
RAM[16'h6327] = 8'h00;
RAM[16'h6328] = 8'h00;
RAM[16'h6329] = 8'h00;
RAM[16'h632A] = 8'h00;
RAM[16'h632B] = 8'h00;
RAM[16'h632C] = 8'h00;
RAM[16'h632D] = 8'h00;
RAM[16'h632E] = 8'h00;
RAM[16'h632F] = 8'h00;
RAM[16'h6330] = 8'h00;
RAM[16'h6331] = 8'h00;
RAM[16'h6332] = 8'h00;
RAM[16'h6333] = 8'h00;
RAM[16'h6334] = 8'h00;
RAM[16'h6335] = 8'h00;
RAM[16'h6336] = 8'h00;
RAM[16'h6337] = 8'h00;
RAM[16'h6338] = 8'h00;
RAM[16'h6339] = 8'h00;
RAM[16'h633A] = 8'h00;
RAM[16'h633B] = 8'h00;
RAM[16'h633C] = 8'h00;
RAM[16'h633D] = 8'h00;
RAM[16'h633E] = 8'h00;
RAM[16'h633F] = 8'h00;
RAM[16'h6340] = 8'h00;
RAM[16'h6341] = 8'h00;
RAM[16'h6342] = 8'h00;
RAM[16'h6343] = 8'h00;
RAM[16'h6344] = 8'h00;
RAM[16'h6345] = 8'h00;
RAM[16'h6346] = 8'h00;
RAM[16'h6347] = 8'h00;
RAM[16'h6348] = 8'h00;
RAM[16'h6349] = 8'h00;
RAM[16'h634A] = 8'h00;
RAM[16'h634B] = 8'h00;
RAM[16'h634C] = 8'h00;
RAM[16'h634D] = 8'h00;
RAM[16'h634E] = 8'h00;
RAM[16'h634F] = 8'h00;
RAM[16'h6350] = 8'h00;
RAM[16'h6351] = 8'h00;
RAM[16'h6352] = 8'h00;
RAM[16'h6353] = 8'h00;
RAM[16'h6354] = 8'h00;
RAM[16'h6355] = 8'h00;
RAM[16'h6356] = 8'h00;
RAM[16'h6357] = 8'h00;
RAM[16'h6358] = 8'h00;
RAM[16'h6359] = 8'h00;
RAM[16'h635A] = 8'h00;
RAM[16'h635B] = 8'h00;
RAM[16'h635C] = 8'h00;
RAM[16'h635D] = 8'h00;
RAM[16'h635E] = 8'h00;
RAM[16'h635F] = 8'h00;
RAM[16'h6360] = 8'h00;
RAM[16'h6361] = 8'h00;
RAM[16'h6362] = 8'h00;
RAM[16'h6363] = 8'h00;
RAM[16'h6364] = 8'h00;
RAM[16'h6365] = 8'h00;
RAM[16'h6366] = 8'h00;
RAM[16'h6367] = 8'h00;
RAM[16'h6368] = 8'h00;
RAM[16'h6369] = 8'h00;
RAM[16'h636A] = 8'h00;
RAM[16'h636B] = 8'h00;
RAM[16'h636C] = 8'h00;
RAM[16'h636D] = 8'h00;
RAM[16'h636E] = 8'h00;
RAM[16'h636F] = 8'h00;
RAM[16'h6370] = 8'h00;
RAM[16'h6371] = 8'h00;
RAM[16'h6372] = 8'h00;
RAM[16'h6373] = 8'h00;
RAM[16'h6374] = 8'h00;
RAM[16'h6375] = 8'h00;
RAM[16'h6376] = 8'h00;
RAM[16'h6377] = 8'h00;
RAM[16'h6378] = 8'h00;
RAM[16'h6379] = 8'h00;
RAM[16'h637A] = 8'h00;
RAM[16'h637B] = 8'h00;
RAM[16'h637C] = 8'h00;
RAM[16'h637D] = 8'h00;
RAM[16'h637E] = 8'h00;
RAM[16'h637F] = 8'h00;
RAM[16'h6380] = 8'h00;
RAM[16'h6381] = 8'h00;
RAM[16'h6382] = 8'h00;
RAM[16'h6383] = 8'h00;
RAM[16'h6384] = 8'h00;
RAM[16'h6385] = 8'h00;
RAM[16'h6386] = 8'h00;
RAM[16'h6387] = 8'h00;
RAM[16'h6388] = 8'h00;
RAM[16'h6389] = 8'h00;
RAM[16'h638A] = 8'h00;
RAM[16'h638B] = 8'h00;
RAM[16'h638C] = 8'h00;
RAM[16'h638D] = 8'h00;
RAM[16'h638E] = 8'h00;
RAM[16'h638F] = 8'h00;
RAM[16'h6390] = 8'h00;
RAM[16'h6391] = 8'h00;
RAM[16'h6392] = 8'h00;
RAM[16'h6393] = 8'h00;
RAM[16'h6394] = 8'h00;
RAM[16'h6395] = 8'h00;
RAM[16'h6396] = 8'h00;
RAM[16'h6397] = 8'h00;
RAM[16'h6398] = 8'h00;
RAM[16'h6399] = 8'h00;
RAM[16'h639A] = 8'h00;
RAM[16'h639B] = 8'h00;
RAM[16'h639C] = 8'h00;
RAM[16'h639D] = 8'h00;
RAM[16'h639E] = 8'h00;
RAM[16'h639F] = 8'h00;
RAM[16'h63A0] = 8'h00;
RAM[16'h63A1] = 8'h00;
RAM[16'h63A2] = 8'h00;
RAM[16'h63A3] = 8'h00;
RAM[16'h63A4] = 8'h00;
RAM[16'h63A5] = 8'h00;
RAM[16'h63A6] = 8'h00;
RAM[16'h63A7] = 8'h00;
RAM[16'h63A8] = 8'h00;
RAM[16'h63A9] = 8'h00;
RAM[16'h63AA] = 8'h00;
RAM[16'h63AB] = 8'h00;
RAM[16'h63AC] = 8'h00;
RAM[16'h63AD] = 8'h00;
RAM[16'h63AE] = 8'h00;
RAM[16'h63AF] = 8'h00;
RAM[16'h63B0] = 8'h00;
RAM[16'h63B1] = 8'h00;
RAM[16'h63B2] = 8'h00;
RAM[16'h63B3] = 8'h00;
RAM[16'h63B4] = 8'h00;
RAM[16'h63B5] = 8'h00;
RAM[16'h63B6] = 8'h00;
RAM[16'h63B7] = 8'h00;
RAM[16'h63B8] = 8'h00;
RAM[16'h63B9] = 8'h00;
RAM[16'h63BA] = 8'h00;
RAM[16'h63BB] = 8'h00;
RAM[16'h63BC] = 8'h00;
RAM[16'h63BD] = 8'h00;
RAM[16'h63BE] = 8'h00;
RAM[16'h63BF] = 8'h00;
RAM[16'h63C0] = 8'h00;
RAM[16'h63C1] = 8'h00;
RAM[16'h63C2] = 8'h00;
RAM[16'h63C3] = 8'h00;
RAM[16'h63C4] = 8'h00;
RAM[16'h63C5] = 8'h00;
RAM[16'h63C6] = 8'h00;
RAM[16'h63C7] = 8'h00;
RAM[16'h63C8] = 8'h00;
RAM[16'h63C9] = 8'h00;
RAM[16'h63CA] = 8'h00;
RAM[16'h63CB] = 8'h00;
RAM[16'h63CC] = 8'h00;
RAM[16'h63CD] = 8'h00;
RAM[16'h63CE] = 8'h00;
RAM[16'h63CF] = 8'h00;
RAM[16'h63D0] = 8'h00;
RAM[16'h63D1] = 8'h00;
RAM[16'h63D2] = 8'h00;
RAM[16'h63D3] = 8'h00;
RAM[16'h63D4] = 8'h00;
RAM[16'h63D5] = 8'h00;
RAM[16'h63D6] = 8'h00;
RAM[16'h63D7] = 8'h00;
RAM[16'h63D8] = 8'h00;
RAM[16'h63D9] = 8'h00;
RAM[16'h63DA] = 8'h00;
RAM[16'h63DB] = 8'h00;
RAM[16'h63DC] = 8'h00;
RAM[16'h63DD] = 8'h00;
RAM[16'h63DE] = 8'h00;
RAM[16'h63DF] = 8'h00;
RAM[16'h63E0] = 8'h00;
RAM[16'h63E1] = 8'h00;
RAM[16'h63E2] = 8'h00;
RAM[16'h63E3] = 8'h00;
RAM[16'h63E4] = 8'h00;
RAM[16'h63E5] = 8'h00;
RAM[16'h63E6] = 8'h00;
RAM[16'h63E7] = 8'h00;
RAM[16'h63E8] = 8'h00;
RAM[16'h63E9] = 8'h00;
RAM[16'h63EA] = 8'h00;
RAM[16'h63EB] = 8'h00;
RAM[16'h63EC] = 8'h00;
RAM[16'h63ED] = 8'h00;
RAM[16'h63EE] = 8'h00;
RAM[16'h63EF] = 8'h00;
RAM[16'h63F0] = 8'h00;
RAM[16'h63F1] = 8'h00;
RAM[16'h63F2] = 8'h00;
RAM[16'h63F3] = 8'h00;
RAM[16'h63F4] = 8'h00;
RAM[16'h63F5] = 8'h00;
RAM[16'h63F6] = 8'h00;
RAM[16'h63F7] = 8'h00;
RAM[16'h63F8] = 8'h00;
RAM[16'h63F9] = 8'h00;
RAM[16'h63FA] = 8'h00;
RAM[16'h63FB] = 8'h00;
RAM[16'h63FC] = 8'h00;
RAM[16'h63FD] = 8'h00;
RAM[16'h63FE] = 8'h00;
RAM[16'h63FF] = 8'h00;
RAM[16'h6400] = 8'h00;
RAM[16'h6401] = 8'h00;
RAM[16'h6402] = 8'h00;
RAM[16'h6403] = 8'h00;
RAM[16'h6404] = 8'h00;
RAM[16'h6405] = 8'h00;
RAM[16'h6406] = 8'h00;
RAM[16'h6407] = 8'h00;
RAM[16'h6408] = 8'h00;
RAM[16'h6409] = 8'h00;
RAM[16'h640A] = 8'h00;
RAM[16'h640B] = 8'h00;
RAM[16'h640C] = 8'h00;
RAM[16'h640D] = 8'h00;
RAM[16'h640E] = 8'h00;
RAM[16'h640F] = 8'h00;
RAM[16'h6410] = 8'h00;
RAM[16'h6411] = 8'h00;
RAM[16'h6412] = 8'h00;
RAM[16'h6413] = 8'h00;
RAM[16'h6414] = 8'h00;
RAM[16'h6415] = 8'h00;
RAM[16'h6416] = 8'h00;
RAM[16'h6417] = 8'h00;
RAM[16'h6418] = 8'h00;
RAM[16'h6419] = 8'h00;
RAM[16'h641A] = 8'h00;
RAM[16'h641B] = 8'h00;
RAM[16'h641C] = 8'h00;
RAM[16'h641D] = 8'h00;
RAM[16'h641E] = 8'h00;
RAM[16'h641F] = 8'h00;
RAM[16'h6420] = 8'h00;
RAM[16'h6421] = 8'h00;
RAM[16'h6422] = 8'h00;
RAM[16'h6423] = 8'h00;
RAM[16'h6424] = 8'h00;
RAM[16'h6425] = 8'h00;
RAM[16'h6426] = 8'h00;
RAM[16'h6427] = 8'h00;
RAM[16'h6428] = 8'h00;
RAM[16'h6429] = 8'h00;
RAM[16'h642A] = 8'h00;
RAM[16'h642B] = 8'h00;
RAM[16'h642C] = 8'h00;
RAM[16'h642D] = 8'h00;
RAM[16'h642E] = 8'h00;
RAM[16'h642F] = 8'h00;
RAM[16'h6430] = 8'h00;
RAM[16'h6431] = 8'h00;
RAM[16'h6432] = 8'h00;
RAM[16'h6433] = 8'h00;
RAM[16'h6434] = 8'h00;
RAM[16'h6435] = 8'h00;
RAM[16'h6436] = 8'h00;
RAM[16'h6437] = 8'h00;
RAM[16'h6438] = 8'h00;
RAM[16'h6439] = 8'h00;
RAM[16'h643A] = 8'h00;
RAM[16'h643B] = 8'h00;
RAM[16'h643C] = 8'h00;
RAM[16'h643D] = 8'h00;
RAM[16'h643E] = 8'h00;
RAM[16'h643F] = 8'h00;
RAM[16'h6440] = 8'h00;
RAM[16'h6441] = 8'h00;
RAM[16'h6442] = 8'h00;
RAM[16'h6443] = 8'h00;
RAM[16'h6444] = 8'h00;
RAM[16'h6445] = 8'h00;
RAM[16'h6446] = 8'h00;
RAM[16'h6447] = 8'h00;
RAM[16'h6448] = 8'h00;
RAM[16'h6449] = 8'h00;
RAM[16'h644A] = 8'h00;
RAM[16'h644B] = 8'h00;
RAM[16'h644C] = 8'h00;
RAM[16'h644D] = 8'h00;
RAM[16'h644E] = 8'h00;
RAM[16'h644F] = 8'h00;
RAM[16'h6450] = 8'h00;
RAM[16'h6451] = 8'h00;
RAM[16'h6452] = 8'h00;
RAM[16'h6453] = 8'h00;
RAM[16'h6454] = 8'h00;
RAM[16'h6455] = 8'h00;
RAM[16'h6456] = 8'h00;
RAM[16'h6457] = 8'h00;
RAM[16'h6458] = 8'h00;
RAM[16'h6459] = 8'h00;
RAM[16'h645A] = 8'h00;
RAM[16'h645B] = 8'h00;
RAM[16'h645C] = 8'h00;
RAM[16'h645D] = 8'h00;
RAM[16'h645E] = 8'h00;
RAM[16'h645F] = 8'h00;
RAM[16'h6460] = 8'h00;
RAM[16'h6461] = 8'h00;
RAM[16'h6462] = 8'h00;
RAM[16'h6463] = 8'h00;
RAM[16'h6464] = 8'h00;
RAM[16'h6465] = 8'h00;
RAM[16'h6466] = 8'h00;
RAM[16'h6467] = 8'h00;
RAM[16'h6468] = 8'h00;
RAM[16'h6469] = 8'h00;
RAM[16'h646A] = 8'h00;
RAM[16'h646B] = 8'h00;
RAM[16'h646C] = 8'h00;
RAM[16'h646D] = 8'h00;
RAM[16'h646E] = 8'h00;
RAM[16'h646F] = 8'h00;
RAM[16'h6470] = 8'h00;
RAM[16'h6471] = 8'h00;
RAM[16'h6472] = 8'h00;
RAM[16'h6473] = 8'h00;
RAM[16'h6474] = 8'h00;
RAM[16'h6475] = 8'h00;
RAM[16'h6476] = 8'h00;
RAM[16'h6477] = 8'h00;
RAM[16'h6478] = 8'h00;
RAM[16'h6479] = 8'h00;
RAM[16'h647A] = 8'h00;
RAM[16'h647B] = 8'h00;
RAM[16'h647C] = 8'h00;
RAM[16'h647D] = 8'h00;
RAM[16'h647E] = 8'h00;
RAM[16'h647F] = 8'h00;
RAM[16'h6480] = 8'h00;
RAM[16'h6481] = 8'h00;
RAM[16'h6482] = 8'h00;
RAM[16'h6483] = 8'h00;
RAM[16'h6484] = 8'h00;
RAM[16'h6485] = 8'h00;
RAM[16'h6486] = 8'h00;
RAM[16'h6487] = 8'h00;
RAM[16'h6488] = 8'h00;
RAM[16'h6489] = 8'h00;
RAM[16'h648A] = 8'h00;
RAM[16'h648B] = 8'h00;
RAM[16'h648C] = 8'h00;
RAM[16'h648D] = 8'h00;
RAM[16'h648E] = 8'h00;
RAM[16'h648F] = 8'h00;
RAM[16'h6490] = 8'h00;
RAM[16'h6491] = 8'h00;
RAM[16'h6492] = 8'h00;
RAM[16'h6493] = 8'h00;
RAM[16'h6494] = 8'h00;
RAM[16'h6495] = 8'h00;
RAM[16'h6496] = 8'h00;
RAM[16'h6497] = 8'h00;
RAM[16'h6498] = 8'h00;
RAM[16'h6499] = 8'h00;
RAM[16'h649A] = 8'h00;
RAM[16'h649B] = 8'h00;
RAM[16'h649C] = 8'h00;
RAM[16'h649D] = 8'h00;
RAM[16'h649E] = 8'h00;
RAM[16'h649F] = 8'h00;
RAM[16'h64A0] = 8'h00;
RAM[16'h64A1] = 8'h00;
RAM[16'h64A2] = 8'h00;
RAM[16'h64A3] = 8'h00;
RAM[16'h64A4] = 8'h00;
RAM[16'h64A5] = 8'h00;
RAM[16'h64A6] = 8'h00;
RAM[16'h64A7] = 8'h00;
RAM[16'h64A8] = 8'h00;
RAM[16'h64A9] = 8'h00;
RAM[16'h64AA] = 8'h00;
RAM[16'h64AB] = 8'h00;
RAM[16'h64AC] = 8'h00;
RAM[16'h64AD] = 8'h00;
RAM[16'h64AE] = 8'h00;
RAM[16'h64AF] = 8'h00;
RAM[16'h64B0] = 8'h00;
RAM[16'h64B1] = 8'h00;
RAM[16'h64B2] = 8'h00;
RAM[16'h64B3] = 8'h00;
RAM[16'h64B4] = 8'h00;
RAM[16'h64B5] = 8'h00;
RAM[16'h64B6] = 8'h00;
RAM[16'h64B7] = 8'h00;
RAM[16'h64B8] = 8'h00;
RAM[16'h64B9] = 8'h00;
RAM[16'h64BA] = 8'h00;
RAM[16'h64BB] = 8'h00;
RAM[16'h64BC] = 8'h00;
RAM[16'h64BD] = 8'h00;
RAM[16'h64BE] = 8'h00;
RAM[16'h64BF] = 8'h00;
RAM[16'h64C0] = 8'h00;
RAM[16'h64C1] = 8'h00;
RAM[16'h64C2] = 8'h00;
RAM[16'h64C3] = 8'h00;
RAM[16'h64C4] = 8'h00;
RAM[16'h64C5] = 8'h00;
RAM[16'h64C6] = 8'h00;
RAM[16'h64C7] = 8'h00;
RAM[16'h64C8] = 8'h00;
RAM[16'h64C9] = 8'h00;
RAM[16'h64CA] = 8'h00;
RAM[16'h64CB] = 8'h00;
RAM[16'h64CC] = 8'h00;
RAM[16'h64CD] = 8'h00;
RAM[16'h64CE] = 8'h00;
RAM[16'h64CF] = 8'h00;
RAM[16'h64D0] = 8'h00;
RAM[16'h64D1] = 8'h00;
RAM[16'h64D2] = 8'h00;
RAM[16'h64D3] = 8'h00;
RAM[16'h64D4] = 8'h00;
RAM[16'h64D5] = 8'h00;
RAM[16'h64D6] = 8'h00;
RAM[16'h64D7] = 8'h00;
RAM[16'h64D8] = 8'h00;
RAM[16'h64D9] = 8'h00;
RAM[16'h64DA] = 8'h00;
RAM[16'h64DB] = 8'h00;
RAM[16'h64DC] = 8'h00;
RAM[16'h64DD] = 8'h00;
RAM[16'h64DE] = 8'h00;
RAM[16'h64DF] = 8'h00;
RAM[16'h64E0] = 8'h00;
RAM[16'h64E1] = 8'h00;
RAM[16'h64E2] = 8'h00;
RAM[16'h64E3] = 8'h00;
RAM[16'h64E4] = 8'h00;
RAM[16'h64E5] = 8'h00;
RAM[16'h64E6] = 8'h00;
RAM[16'h64E7] = 8'h00;
RAM[16'h64E8] = 8'h00;
RAM[16'h64E9] = 8'h00;
RAM[16'h64EA] = 8'h00;
RAM[16'h64EB] = 8'h00;
RAM[16'h64EC] = 8'h00;
RAM[16'h64ED] = 8'h00;
RAM[16'h64EE] = 8'h00;
RAM[16'h64EF] = 8'h00;
RAM[16'h64F0] = 8'h00;
RAM[16'h64F1] = 8'h00;
RAM[16'h64F2] = 8'h00;
RAM[16'h64F3] = 8'h00;
RAM[16'h64F4] = 8'h00;
RAM[16'h64F5] = 8'h00;
RAM[16'h64F6] = 8'h00;
RAM[16'h64F7] = 8'h00;
RAM[16'h64F8] = 8'h00;
RAM[16'h64F9] = 8'h00;
RAM[16'h64FA] = 8'h00;
RAM[16'h64FB] = 8'h00;
RAM[16'h64FC] = 8'h00;
RAM[16'h64FD] = 8'h00;
RAM[16'h64FE] = 8'h00;
RAM[16'h64FF] = 8'h00;
RAM[16'h6500] = 8'h00;
RAM[16'h6501] = 8'h00;
RAM[16'h6502] = 8'h00;
RAM[16'h6503] = 8'h00;
RAM[16'h6504] = 8'h00;
RAM[16'h6505] = 8'h00;
RAM[16'h6506] = 8'h00;
RAM[16'h6507] = 8'h00;
RAM[16'h6508] = 8'h00;
RAM[16'h6509] = 8'h00;
RAM[16'h650A] = 8'h00;
RAM[16'h650B] = 8'h00;
RAM[16'h650C] = 8'h00;
RAM[16'h650D] = 8'h00;
RAM[16'h650E] = 8'h00;
RAM[16'h650F] = 8'h00;
RAM[16'h6510] = 8'h00;
RAM[16'h6511] = 8'h00;
RAM[16'h6512] = 8'h00;
RAM[16'h6513] = 8'h00;
RAM[16'h6514] = 8'h00;
RAM[16'h6515] = 8'h00;
RAM[16'h6516] = 8'h00;
RAM[16'h6517] = 8'h00;
RAM[16'h6518] = 8'h00;
RAM[16'h6519] = 8'h00;
RAM[16'h651A] = 8'h00;
RAM[16'h651B] = 8'h00;
RAM[16'h651C] = 8'h00;
RAM[16'h651D] = 8'h00;
RAM[16'h651E] = 8'h00;
RAM[16'h651F] = 8'h00;
RAM[16'h6520] = 8'h00;
RAM[16'h6521] = 8'h00;
RAM[16'h6522] = 8'h00;
RAM[16'h6523] = 8'h00;
RAM[16'h6524] = 8'h00;
RAM[16'h6525] = 8'h00;
RAM[16'h6526] = 8'h00;
RAM[16'h6527] = 8'h00;
RAM[16'h6528] = 8'h00;
RAM[16'h6529] = 8'h00;
RAM[16'h652A] = 8'h00;
RAM[16'h652B] = 8'h00;
RAM[16'h652C] = 8'h00;
RAM[16'h652D] = 8'h00;
RAM[16'h652E] = 8'h00;
RAM[16'h652F] = 8'h00;
RAM[16'h6530] = 8'h00;
RAM[16'h6531] = 8'h00;
RAM[16'h6532] = 8'h00;
RAM[16'h6533] = 8'h00;
RAM[16'h6534] = 8'h00;
RAM[16'h6535] = 8'h00;
RAM[16'h6536] = 8'h00;
RAM[16'h6537] = 8'h00;
RAM[16'h6538] = 8'h00;
RAM[16'h6539] = 8'h00;
RAM[16'h653A] = 8'h00;
RAM[16'h653B] = 8'h00;
RAM[16'h653C] = 8'h00;
RAM[16'h653D] = 8'h00;
RAM[16'h653E] = 8'h00;
RAM[16'h653F] = 8'h00;
RAM[16'h6540] = 8'h00;
RAM[16'h6541] = 8'h00;
RAM[16'h6542] = 8'h00;
RAM[16'h6543] = 8'h00;
RAM[16'h6544] = 8'h00;
RAM[16'h6545] = 8'h00;
RAM[16'h6546] = 8'h00;
RAM[16'h6547] = 8'h00;
RAM[16'h6548] = 8'h00;
RAM[16'h6549] = 8'h00;
RAM[16'h654A] = 8'h00;
RAM[16'h654B] = 8'h00;
RAM[16'h654C] = 8'h00;
RAM[16'h654D] = 8'h00;
RAM[16'h654E] = 8'h00;
RAM[16'h654F] = 8'h00;
RAM[16'h6550] = 8'h00;
RAM[16'h6551] = 8'h00;
RAM[16'h6552] = 8'h00;
RAM[16'h6553] = 8'h00;
RAM[16'h6554] = 8'h00;
RAM[16'h6555] = 8'h00;
RAM[16'h6556] = 8'h00;
RAM[16'h6557] = 8'h00;
RAM[16'h6558] = 8'h00;
RAM[16'h6559] = 8'h00;
RAM[16'h655A] = 8'h00;
RAM[16'h655B] = 8'h00;
RAM[16'h655C] = 8'h00;
RAM[16'h655D] = 8'h00;
RAM[16'h655E] = 8'h00;
RAM[16'h655F] = 8'h00;
RAM[16'h6560] = 8'h00;
RAM[16'h6561] = 8'h00;
RAM[16'h6562] = 8'h00;
RAM[16'h6563] = 8'h00;
RAM[16'h6564] = 8'h00;
RAM[16'h6565] = 8'h00;
RAM[16'h6566] = 8'h00;
RAM[16'h6567] = 8'h00;
RAM[16'h6568] = 8'h00;
RAM[16'h6569] = 8'h00;
RAM[16'h656A] = 8'h00;
RAM[16'h656B] = 8'h00;
RAM[16'h656C] = 8'h00;
RAM[16'h656D] = 8'h00;
RAM[16'h656E] = 8'h00;
RAM[16'h656F] = 8'h00;
RAM[16'h6570] = 8'h00;
RAM[16'h6571] = 8'h00;
RAM[16'h6572] = 8'h00;
RAM[16'h6573] = 8'h00;
RAM[16'h6574] = 8'h00;
RAM[16'h6575] = 8'h00;
RAM[16'h6576] = 8'h00;
RAM[16'h6577] = 8'h00;
RAM[16'h6578] = 8'h00;
RAM[16'h6579] = 8'h00;
RAM[16'h657A] = 8'h00;
RAM[16'h657B] = 8'h00;
RAM[16'h657C] = 8'h00;
RAM[16'h657D] = 8'h00;
RAM[16'h657E] = 8'h00;
RAM[16'h657F] = 8'h00;
RAM[16'h6580] = 8'h00;
RAM[16'h6581] = 8'h00;
RAM[16'h6582] = 8'h00;
RAM[16'h6583] = 8'h00;
RAM[16'h6584] = 8'h00;
RAM[16'h6585] = 8'h00;
RAM[16'h6586] = 8'h00;
RAM[16'h6587] = 8'h00;
RAM[16'h6588] = 8'h00;
RAM[16'h6589] = 8'h00;
RAM[16'h658A] = 8'h00;
RAM[16'h658B] = 8'h00;
RAM[16'h658C] = 8'h00;
RAM[16'h658D] = 8'h00;
RAM[16'h658E] = 8'h00;
RAM[16'h658F] = 8'h00;
RAM[16'h6590] = 8'h00;
RAM[16'h6591] = 8'h00;
RAM[16'h6592] = 8'h00;
RAM[16'h6593] = 8'h00;
RAM[16'h6594] = 8'h00;
RAM[16'h6595] = 8'h00;
RAM[16'h6596] = 8'h00;
RAM[16'h6597] = 8'h00;
RAM[16'h6598] = 8'h00;
RAM[16'h6599] = 8'h00;
RAM[16'h659A] = 8'h00;
RAM[16'h659B] = 8'h00;
RAM[16'h659C] = 8'h00;
RAM[16'h659D] = 8'h00;
RAM[16'h659E] = 8'h00;
RAM[16'h659F] = 8'h00;
RAM[16'h65A0] = 8'h00;
RAM[16'h65A1] = 8'h00;
RAM[16'h65A2] = 8'h00;
RAM[16'h65A3] = 8'h00;
RAM[16'h65A4] = 8'h00;
RAM[16'h65A5] = 8'h00;
RAM[16'h65A6] = 8'h00;
RAM[16'h65A7] = 8'h00;
RAM[16'h65A8] = 8'h00;
RAM[16'h65A9] = 8'h00;
RAM[16'h65AA] = 8'h00;
RAM[16'h65AB] = 8'h00;
RAM[16'h65AC] = 8'h00;
RAM[16'h65AD] = 8'h00;
RAM[16'h65AE] = 8'h00;
RAM[16'h65AF] = 8'h00;
RAM[16'h65B0] = 8'h00;
RAM[16'h65B1] = 8'h00;
RAM[16'h65B2] = 8'h00;
RAM[16'h65B3] = 8'h00;
RAM[16'h65B4] = 8'h00;
RAM[16'h65B5] = 8'h00;
RAM[16'h65B6] = 8'h00;
RAM[16'h65B7] = 8'h00;
RAM[16'h65B8] = 8'h00;
RAM[16'h65B9] = 8'h00;
RAM[16'h65BA] = 8'h00;
RAM[16'h65BB] = 8'h00;
RAM[16'h65BC] = 8'h00;
RAM[16'h65BD] = 8'h00;
RAM[16'h65BE] = 8'h00;
RAM[16'h65BF] = 8'h00;
RAM[16'h65C0] = 8'h00;
RAM[16'h65C1] = 8'h00;
RAM[16'h65C2] = 8'h00;
RAM[16'h65C3] = 8'h00;
RAM[16'h65C4] = 8'h00;
RAM[16'h65C5] = 8'h00;
RAM[16'h65C6] = 8'h00;
RAM[16'h65C7] = 8'h00;
RAM[16'h65C8] = 8'h00;
RAM[16'h65C9] = 8'h00;
RAM[16'h65CA] = 8'h00;
RAM[16'h65CB] = 8'h00;
RAM[16'h65CC] = 8'h00;
RAM[16'h65CD] = 8'h00;
RAM[16'h65CE] = 8'h00;
RAM[16'h65CF] = 8'h00;
RAM[16'h65D0] = 8'h00;
RAM[16'h65D1] = 8'h00;
RAM[16'h65D2] = 8'h00;
RAM[16'h65D3] = 8'h00;
RAM[16'h65D4] = 8'h00;
RAM[16'h65D5] = 8'h00;
RAM[16'h65D6] = 8'h00;
RAM[16'h65D7] = 8'h00;
RAM[16'h65D8] = 8'h00;
RAM[16'h65D9] = 8'h00;
RAM[16'h65DA] = 8'h00;
RAM[16'h65DB] = 8'h00;
RAM[16'h65DC] = 8'h00;
RAM[16'h65DD] = 8'h00;
RAM[16'h65DE] = 8'h00;
RAM[16'h65DF] = 8'h00;
RAM[16'h65E0] = 8'h00;
RAM[16'h65E1] = 8'h00;
RAM[16'h65E2] = 8'h00;
RAM[16'h65E3] = 8'h00;
RAM[16'h65E4] = 8'h00;
RAM[16'h65E5] = 8'h00;
RAM[16'h65E6] = 8'h00;
RAM[16'h65E7] = 8'h00;
RAM[16'h65E8] = 8'h00;
RAM[16'h65E9] = 8'h00;
RAM[16'h65EA] = 8'h00;
RAM[16'h65EB] = 8'h00;
RAM[16'h65EC] = 8'h00;
RAM[16'h65ED] = 8'h00;
RAM[16'h65EE] = 8'h00;
RAM[16'h65EF] = 8'h00;
RAM[16'h65F0] = 8'h00;
RAM[16'h65F1] = 8'h00;
RAM[16'h65F2] = 8'h00;
RAM[16'h65F3] = 8'h00;
RAM[16'h65F4] = 8'h00;
RAM[16'h65F5] = 8'h00;
RAM[16'h65F6] = 8'h00;
RAM[16'h65F7] = 8'h00;
RAM[16'h65F8] = 8'h00;
RAM[16'h65F9] = 8'h00;
RAM[16'h65FA] = 8'h00;
RAM[16'h65FB] = 8'h00;
RAM[16'h65FC] = 8'h00;
RAM[16'h65FD] = 8'h00;
RAM[16'h65FE] = 8'h00;
RAM[16'h65FF] = 8'h00;
RAM[16'h6600] = 8'h00;
RAM[16'h6601] = 8'h00;
RAM[16'h6602] = 8'h00;
RAM[16'h6603] = 8'h00;
RAM[16'h6604] = 8'h00;
RAM[16'h6605] = 8'h00;
RAM[16'h6606] = 8'h00;
RAM[16'h6607] = 8'h00;
RAM[16'h6608] = 8'h00;
RAM[16'h6609] = 8'h00;
RAM[16'h660A] = 8'h00;
RAM[16'h660B] = 8'h00;
RAM[16'h660C] = 8'h00;
RAM[16'h660D] = 8'h00;
RAM[16'h660E] = 8'h00;
RAM[16'h660F] = 8'h00;
RAM[16'h6610] = 8'h00;
RAM[16'h6611] = 8'h00;
RAM[16'h6612] = 8'h00;
RAM[16'h6613] = 8'h00;
RAM[16'h6614] = 8'h00;
RAM[16'h6615] = 8'h00;
RAM[16'h6616] = 8'h00;
RAM[16'h6617] = 8'h00;
RAM[16'h6618] = 8'h00;
RAM[16'h6619] = 8'h00;
RAM[16'h661A] = 8'h00;
RAM[16'h661B] = 8'h00;
RAM[16'h661C] = 8'h00;
RAM[16'h661D] = 8'h00;
RAM[16'h661E] = 8'h00;
RAM[16'h661F] = 8'h00;
RAM[16'h6620] = 8'h00;
RAM[16'h6621] = 8'h00;
RAM[16'h6622] = 8'h00;
RAM[16'h6623] = 8'h00;
RAM[16'h6624] = 8'h00;
RAM[16'h6625] = 8'h00;
RAM[16'h6626] = 8'h00;
RAM[16'h6627] = 8'h00;
RAM[16'h6628] = 8'h00;
RAM[16'h6629] = 8'h00;
RAM[16'h662A] = 8'h00;
RAM[16'h662B] = 8'h00;
RAM[16'h662C] = 8'h00;
RAM[16'h662D] = 8'h00;
RAM[16'h662E] = 8'h00;
RAM[16'h662F] = 8'h00;
RAM[16'h6630] = 8'h00;
RAM[16'h6631] = 8'h00;
RAM[16'h6632] = 8'h00;
RAM[16'h6633] = 8'h00;
RAM[16'h6634] = 8'h00;
RAM[16'h6635] = 8'h00;
RAM[16'h6636] = 8'h00;
RAM[16'h6637] = 8'h00;
RAM[16'h6638] = 8'h00;
RAM[16'h6639] = 8'h00;
RAM[16'h663A] = 8'h00;
RAM[16'h663B] = 8'h00;
RAM[16'h663C] = 8'h00;
RAM[16'h663D] = 8'h00;
RAM[16'h663E] = 8'h00;
RAM[16'h663F] = 8'h00;
RAM[16'h6640] = 8'h00;
RAM[16'h6641] = 8'h00;
RAM[16'h6642] = 8'h00;
RAM[16'h6643] = 8'h00;
RAM[16'h6644] = 8'h00;
RAM[16'h6645] = 8'h00;
RAM[16'h6646] = 8'h00;
RAM[16'h6647] = 8'h00;
RAM[16'h6648] = 8'h00;
RAM[16'h6649] = 8'h00;
RAM[16'h664A] = 8'h00;
RAM[16'h664B] = 8'h00;
RAM[16'h664C] = 8'h00;
RAM[16'h664D] = 8'h00;
RAM[16'h664E] = 8'h00;
RAM[16'h664F] = 8'h00;
RAM[16'h6650] = 8'h00;
RAM[16'h6651] = 8'h00;
RAM[16'h6652] = 8'h00;
RAM[16'h6653] = 8'h00;
RAM[16'h6654] = 8'h00;
RAM[16'h6655] = 8'h00;
RAM[16'h6656] = 8'h00;
RAM[16'h6657] = 8'h00;
RAM[16'h6658] = 8'h00;
RAM[16'h6659] = 8'h00;
RAM[16'h665A] = 8'h00;
RAM[16'h665B] = 8'h00;
RAM[16'h665C] = 8'h00;
RAM[16'h665D] = 8'h00;
RAM[16'h665E] = 8'h00;
RAM[16'h665F] = 8'h00;
RAM[16'h6660] = 8'h00;
RAM[16'h6661] = 8'h00;
RAM[16'h6662] = 8'h00;
RAM[16'h6663] = 8'h00;
RAM[16'h6664] = 8'h00;
RAM[16'h6665] = 8'h00;
RAM[16'h6666] = 8'h00;
RAM[16'h6667] = 8'h00;
RAM[16'h6668] = 8'h00;
RAM[16'h6669] = 8'h00;
RAM[16'h666A] = 8'h00;
RAM[16'h666B] = 8'h00;
RAM[16'h666C] = 8'h00;
RAM[16'h666D] = 8'h00;
RAM[16'h666E] = 8'h00;
RAM[16'h666F] = 8'h00;
RAM[16'h6670] = 8'h00;
RAM[16'h6671] = 8'h00;
RAM[16'h6672] = 8'h00;
RAM[16'h6673] = 8'h00;
RAM[16'h6674] = 8'h00;
RAM[16'h6675] = 8'h00;
RAM[16'h6676] = 8'h00;
RAM[16'h6677] = 8'h00;
RAM[16'h6678] = 8'h00;
RAM[16'h6679] = 8'h00;
RAM[16'h667A] = 8'h00;
RAM[16'h667B] = 8'h00;
RAM[16'h667C] = 8'h00;
RAM[16'h667D] = 8'h00;
RAM[16'h667E] = 8'h00;
RAM[16'h667F] = 8'h00;
RAM[16'h6680] = 8'h00;
RAM[16'h6681] = 8'h00;
RAM[16'h6682] = 8'h00;
RAM[16'h6683] = 8'h00;
RAM[16'h6684] = 8'h00;
RAM[16'h6685] = 8'h00;
RAM[16'h6686] = 8'h00;
RAM[16'h6687] = 8'h00;
RAM[16'h6688] = 8'h00;
RAM[16'h6689] = 8'h00;
RAM[16'h668A] = 8'h00;
RAM[16'h668B] = 8'h00;
RAM[16'h668C] = 8'h00;
RAM[16'h668D] = 8'h00;
RAM[16'h668E] = 8'h00;
RAM[16'h668F] = 8'h00;
RAM[16'h6690] = 8'h00;
RAM[16'h6691] = 8'h00;
RAM[16'h6692] = 8'h00;
RAM[16'h6693] = 8'h00;
RAM[16'h6694] = 8'h00;
RAM[16'h6695] = 8'h00;
RAM[16'h6696] = 8'h00;
RAM[16'h6697] = 8'h00;
RAM[16'h6698] = 8'h00;
RAM[16'h6699] = 8'h00;
RAM[16'h669A] = 8'h00;
RAM[16'h669B] = 8'h00;
RAM[16'h669C] = 8'h00;
RAM[16'h669D] = 8'h00;
RAM[16'h669E] = 8'h00;
RAM[16'h669F] = 8'h00;
RAM[16'h66A0] = 8'h00;
RAM[16'h66A1] = 8'h00;
RAM[16'h66A2] = 8'h00;
RAM[16'h66A3] = 8'h00;
RAM[16'h66A4] = 8'h00;
RAM[16'h66A5] = 8'h00;
RAM[16'h66A6] = 8'h00;
RAM[16'h66A7] = 8'h00;
RAM[16'h66A8] = 8'h00;
RAM[16'h66A9] = 8'h00;
RAM[16'h66AA] = 8'h00;
RAM[16'h66AB] = 8'h00;
RAM[16'h66AC] = 8'h00;
RAM[16'h66AD] = 8'h00;
RAM[16'h66AE] = 8'h00;
RAM[16'h66AF] = 8'h00;
RAM[16'h66B0] = 8'h00;
RAM[16'h66B1] = 8'h00;
RAM[16'h66B2] = 8'h00;
RAM[16'h66B3] = 8'h00;
RAM[16'h66B4] = 8'h00;
RAM[16'h66B5] = 8'h00;
RAM[16'h66B6] = 8'h00;
RAM[16'h66B7] = 8'h00;
RAM[16'h66B8] = 8'h00;
RAM[16'h66B9] = 8'h00;
RAM[16'h66BA] = 8'h00;
RAM[16'h66BB] = 8'h00;
RAM[16'h66BC] = 8'h00;
RAM[16'h66BD] = 8'h00;
RAM[16'h66BE] = 8'h00;
RAM[16'h66BF] = 8'h00;
RAM[16'h66C0] = 8'h00;
RAM[16'h66C1] = 8'h00;
RAM[16'h66C2] = 8'h00;
RAM[16'h66C3] = 8'h00;
RAM[16'h66C4] = 8'h00;
RAM[16'h66C5] = 8'h00;
RAM[16'h66C6] = 8'h00;
RAM[16'h66C7] = 8'h00;
RAM[16'h66C8] = 8'h00;
RAM[16'h66C9] = 8'h00;
RAM[16'h66CA] = 8'h00;
RAM[16'h66CB] = 8'h00;
RAM[16'h66CC] = 8'h00;
RAM[16'h66CD] = 8'h00;
RAM[16'h66CE] = 8'h00;
RAM[16'h66CF] = 8'h00;
RAM[16'h66D0] = 8'h00;
RAM[16'h66D1] = 8'h00;
RAM[16'h66D2] = 8'h00;
RAM[16'h66D3] = 8'h00;
RAM[16'h66D4] = 8'h00;
RAM[16'h66D5] = 8'h00;
RAM[16'h66D6] = 8'h00;
RAM[16'h66D7] = 8'h00;
RAM[16'h66D8] = 8'h00;
RAM[16'h66D9] = 8'h00;
RAM[16'h66DA] = 8'h00;
RAM[16'h66DB] = 8'h00;
RAM[16'h66DC] = 8'h00;
RAM[16'h66DD] = 8'h00;
RAM[16'h66DE] = 8'h00;
RAM[16'h66DF] = 8'h00;
RAM[16'h66E0] = 8'h00;
RAM[16'h66E1] = 8'h00;
RAM[16'h66E2] = 8'h00;
RAM[16'h66E3] = 8'h00;
RAM[16'h66E4] = 8'h00;
RAM[16'h66E5] = 8'h00;
RAM[16'h66E6] = 8'h00;
RAM[16'h66E7] = 8'h00;
RAM[16'h66E8] = 8'h00;
RAM[16'h66E9] = 8'h00;
RAM[16'h66EA] = 8'h00;
RAM[16'h66EB] = 8'h00;
RAM[16'h66EC] = 8'h00;
RAM[16'h66ED] = 8'h00;
RAM[16'h66EE] = 8'h00;
RAM[16'h66EF] = 8'h00;
RAM[16'h66F0] = 8'h00;
RAM[16'h66F1] = 8'h00;
RAM[16'h66F2] = 8'h00;
RAM[16'h66F3] = 8'h00;
RAM[16'h66F4] = 8'h00;
RAM[16'h66F5] = 8'h00;
RAM[16'h66F6] = 8'h00;
RAM[16'h66F7] = 8'h00;
RAM[16'h66F8] = 8'h00;
RAM[16'h66F9] = 8'h00;
RAM[16'h66FA] = 8'h00;
RAM[16'h66FB] = 8'h00;
RAM[16'h66FC] = 8'h00;
RAM[16'h66FD] = 8'h00;
RAM[16'h66FE] = 8'h00;
RAM[16'h66FF] = 8'h00;
RAM[16'h6700] = 8'h00;
RAM[16'h6701] = 8'h00;
RAM[16'h6702] = 8'h00;
RAM[16'h6703] = 8'h00;
RAM[16'h6704] = 8'h00;
RAM[16'h6705] = 8'h00;
RAM[16'h6706] = 8'h00;
RAM[16'h6707] = 8'h00;
RAM[16'h6708] = 8'h00;
RAM[16'h6709] = 8'h00;
RAM[16'h670A] = 8'h00;
RAM[16'h670B] = 8'h00;
RAM[16'h670C] = 8'h00;
RAM[16'h670D] = 8'h00;
RAM[16'h670E] = 8'h00;
RAM[16'h670F] = 8'h00;
RAM[16'h6710] = 8'h00;
RAM[16'h6711] = 8'h00;
RAM[16'h6712] = 8'h00;
RAM[16'h6713] = 8'h00;
RAM[16'h6714] = 8'h00;
RAM[16'h6715] = 8'h00;
RAM[16'h6716] = 8'h00;
RAM[16'h6717] = 8'h00;
RAM[16'h6718] = 8'h00;
RAM[16'h6719] = 8'h00;
RAM[16'h671A] = 8'h00;
RAM[16'h671B] = 8'h00;
RAM[16'h671C] = 8'h00;
RAM[16'h671D] = 8'h00;
RAM[16'h671E] = 8'h00;
RAM[16'h671F] = 8'h00;
RAM[16'h6720] = 8'h00;
RAM[16'h6721] = 8'h00;
RAM[16'h6722] = 8'h00;
RAM[16'h6723] = 8'h00;
RAM[16'h6724] = 8'h00;
RAM[16'h6725] = 8'h00;
RAM[16'h6726] = 8'h00;
RAM[16'h6727] = 8'h00;
RAM[16'h6728] = 8'h00;
RAM[16'h6729] = 8'h00;
RAM[16'h672A] = 8'h00;
RAM[16'h672B] = 8'h00;
RAM[16'h672C] = 8'h00;
RAM[16'h672D] = 8'h00;
RAM[16'h672E] = 8'h00;
RAM[16'h672F] = 8'h00;
RAM[16'h6730] = 8'h00;
RAM[16'h6731] = 8'h00;
RAM[16'h6732] = 8'h00;
RAM[16'h6733] = 8'h00;
RAM[16'h6734] = 8'h00;
RAM[16'h6735] = 8'h00;
RAM[16'h6736] = 8'h00;
RAM[16'h6737] = 8'h00;
RAM[16'h6738] = 8'h00;
RAM[16'h6739] = 8'h00;
RAM[16'h673A] = 8'h00;
RAM[16'h673B] = 8'h00;
RAM[16'h673C] = 8'h00;
RAM[16'h673D] = 8'h00;
RAM[16'h673E] = 8'h00;
RAM[16'h673F] = 8'h00;
RAM[16'h6740] = 8'h00;
RAM[16'h6741] = 8'h00;
RAM[16'h6742] = 8'h00;
RAM[16'h6743] = 8'h00;
RAM[16'h6744] = 8'h00;
RAM[16'h6745] = 8'h00;
RAM[16'h6746] = 8'h00;
RAM[16'h6747] = 8'h00;
RAM[16'h6748] = 8'h00;
RAM[16'h6749] = 8'h00;
RAM[16'h674A] = 8'h00;
RAM[16'h674B] = 8'h00;
RAM[16'h674C] = 8'h00;
RAM[16'h674D] = 8'h00;
RAM[16'h674E] = 8'h00;
RAM[16'h674F] = 8'h00;
RAM[16'h6750] = 8'h00;
RAM[16'h6751] = 8'h00;
RAM[16'h6752] = 8'h00;
RAM[16'h6753] = 8'h00;
RAM[16'h6754] = 8'h00;
RAM[16'h6755] = 8'h00;
RAM[16'h6756] = 8'h00;
RAM[16'h6757] = 8'h00;
RAM[16'h6758] = 8'h00;
RAM[16'h6759] = 8'h00;
RAM[16'h675A] = 8'h00;
RAM[16'h675B] = 8'h00;
RAM[16'h675C] = 8'h00;
RAM[16'h675D] = 8'h00;
RAM[16'h675E] = 8'h00;
RAM[16'h675F] = 8'h00;
RAM[16'h6760] = 8'h00;
RAM[16'h6761] = 8'h00;
RAM[16'h6762] = 8'h00;
RAM[16'h6763] = 8'h00;
RAM[16'h6764] = 8'h00;
RAM[16'h6765] = 8'h00;
RAM[16'h6766] = 8'h00;
RAM[16'h6767] = 8'h00;
RAM[16'h6768] = 8'h00;
RAM[16'h6769] = 8'h00;
RAM[16'h676A] = 8'h00;
RAM[16'h676B] = 8'h00;
RAM[16'h676C] = 8'h00;
RAM[16'h676D] = 8'h00;
RAM[16'h676E] = 8'h00;
RAM[16'h676F] = 8'h00;
RAM[16'h6770] = 8'h00;
RAM[16'h6771] = 8'h00;
RAM[16'h6772] = 8'h00;
RAM[16'h6773] = 8'h00;
RAM[16'h6774] = 8'h00;
RAM[16'h6775] = 8'h00;
RAM[16'h6776] = 8'h00;
RAM[16'h6777] = 8'h00;
RAM[16'h6778] = 8'h00;
RAM[16'h6779] = 8'h00;
RAM[16'h677A] = 8'h00;
RAM[16'h677B] = 8'h00;
RAM[16'h677C] = 8'h00;
RAM[16'h677D] = 8'h00;
RAM[16'h677E] = 8'h00;
RAM[16'h677F] = 8'h00;
RAM[16'h6780] = 8'h00;
RAM[16'h6781] = 8'h00;
RAM[16'h6782] = 8'h00;
RAM[16'h6783] = 8'h00;
RAM[16'h6784] = 8'h00;
RAM[16'h6785] = 8'h00;
RAM[16'h6786] = 8'h00;
RAM[16'h6787] = 8'h00;
RAM[16'h6788] = 8'h00;
RAM[16'h6789] = 8'h00;
RAM[16'h678A] = 8'h00;
RAM[16'h678B] = 8'h00;
RAM[16'h678C] = 8'h00;
RAM[16'h678D] = 8'h00;
RAM[16'h678E] = 8'h00;
RAM[16'h678F] = 8'h00;
RAM[16'h6790] = 8'h00;
RAM[16'h6791] = 8'h00;
RAM[16'h6792] = 8'h00;
RAM[16'h6793] = 8'h00;
RAM[16'h6794] = 8'h00;
RAM[16'h6795] = 8'h00;
RAM[16'h6796] = 8'h00;
RAM[16'h6797] = 8'h00;
RAM[16'h6798] = 8'h00;
RAM[16'h6799] = 8'h00;
RAM[16'h679A] = 8'h00;
RAM[16'h679B] = 8'h00;
RAM[16'h679C] = 8'h00;
RAM[16'h679D] = 8'h00;
RAM[16'h679E] = 8'h00;
RAM[16'h679F] = 8'h00;
RAM[16'h67A0] = 8'h00;
RAM[16'h67A1] = 8'h00;
RAM[16'h67A2] = 8'h00;
RAM[16'h67A3] = 8'h00;
RAM[16'h67A4] = 8'h00;
RAM[16'h67A5] = 8'h00;
RAM[16'h67A6] = 8'h00;
RAM[16'h67A7] = 8'h00;
RAM[16'h67A8] = 8'h00;
RAM[16'h67A9] = 8'h00;
RAM[16'h67AA] = 8'h00;
RAM[16'h67AB] = 8'h00;
RAM[16'h67AC] = 8'h00;
RAM[16'h67AD] = 8'h00;
RAM[16'h67AE] = 8'h00;
RAM[16'h67AF] = 8'h00;
RAM[16'h67B0] = 8'h00;
RAM[16'h67B1] = 8'h00;
RAM[16'h67B2] = 8'h00;
RAM[16'h67B3] = 8'h00;
RAM[16'h67B4] = 8'h00;
RAM[16'h67B5] = 8'h00;
RAM[16'h67B6] = 8'h00;
RAM[16'h67B7] = 8'h00;
RAM[16'h67B8] = 8'h00;
RAM[16'h67B9] = 8'h00;
RAM[16'h67BA] = 8'h00;
RAM[16'h67BB] = 8'h00;
RAM[16'h67BC] = 8'h00;
RAM[16'h67BD] = 8'h00;
RAM[16'h67BE] = 8'h00;
RAM[16'h67BF] = 8'h00;
RAM[16'h67C0] = 8'h00;
RAM[16'h67C1] = 8'h00;
RAM[16'h67C2] = 8'h00;
RAM[16'h67C3] = 8'h00;
RAM[16'h67C4] = 8'h00;
RAM[16'h67C5] = 8'h00;
RAM[16'h67C6] = 8'h00;
RAM[16'h67C7] = 8'h00;
RAM[16'h67C8] = 8'h00;
RAM[16'h67C9] = 8'h00;
RAM[16'h67CA] = 8'h00;
RAM[16'h67CB] = 8'h00;
RAM[16'h67CC] = 8'h00;
RAM[16'h67CD] = 8'h00;
RAM[16'h67CE] = 8'h00;
RAM[16'h67CF] = 8'h00;
RAM[16'h67D0] = 8'h00;
RAM[16'h67D1] = 8'h00;
RAM[16'h67D2] = 8'h00;
RAM[16'h67D3] = 8'h00;
RAM[16'h67D4] = 8'h00;
RAM[16'h67D5] = 8'h00;
RAM[16'h67D6] = 8'h00;
RAM[16'h67D7] = 8'h00;
RAM[16'h67D8] = 8'h00;
RAM[16'h67D9] = 8'h00;
RAM[16'h67DA] = 8'h00;
RAM[16'h67DB] = 8'h00;
RAM[16'h67DC] = 8'h00;
RAM[16'h67DD] = 8'h00;
RAM[16'h67DE] = 8'h00;
RAM[16'h67DF] = 8'h00;
RAM[16'h67E0] = 8'h00;
RAM[16'h67E1] = 8'h00;
RAM[16'h67E2] = 8'h00;
RAM[16'h67E3] = 8'h00;
RAM[16'h67E4] = 8'h00;
RAM[16'h67E5] = 8'h00;
RAM[16'h67E6] = 8'h00;
RAM[16'h67E7] = 8'h00;
RAM[16'h67E8] = 8'h00;
RAM[16'h67E9] = 8'h00;
RAM[16'h67EA] = 8'h00;
RAM[16'h67EB] = 8'h00;
RAM[16'h67EC] = 8'h00;
RAM[16'h67ED] = 8'h00;
RAM[16'h67EE] = 8'h00;
RAM[16'h67EF] = 8'h00;
RAM[16'h67F0] = 8'h00;
RAM[16'h67F1] = 8'h00;
RAM[16'h67F2] = 8'h00;
RAM[16'h67F3] = 8'h00;
RAM[16'h67F4] = 8'h00;
RAM[16'h67F5] = 8'h00;
RAM[16'h67F6] = 8'h00;
RAM[16'h67F7] = 8'h00;
RAM[16'h67F8] = 8'h00;
RAM[16'h67F9] = 8'h00;
RAM[16'h67FA] = 8'h00;
RAM[16'h67FB] = 8'h00;
RAM[16'h67FC] = 8'h00;
RAM[16'h67FD] = 8'h00;
RAM[16'h67FE] = 8'h00;
RAM[16'h67FF] = 8'h00;
RAM[16'h6800] = 8'h00;
RAM[16'h6801] = 8'h00;
RAM[16'h6802] = 8'h00;
RAM[16'h6803] = 8'h00;
RAM[16'h6804] = 8'h00;
RAM[16'h6805] = 8'h00;
RAM[16'h6806] = 8'h00;
RAM[16'h6807] = 8'h00;
RAM[16'h6808] = 8'h00;
RAM[16'h6809] = 8'h00;
RAM[16'h680A] = 8'h00;
RAM[16'h680B] = 8'h00;
RAM[16'h680C] = 8'h00;
RAM[16'h680D] = 8'h00;
RAM[16'h680E] = 8'h00;
RAM[16'h680F] = 8'h00;
RAM[16'h6810] = 8'h00;
RAM[16'h6811] = 8'h00;
RAM[16'h6812] = 8'h00;
RAM[16'h6813] = 8'h00;
RAM[16'h6814] = 8'h00;
RAM[16'h6815] = 8'h00;
RAM[16'h6816] = 8'h00;
RAM[16'h6817] = 8'h00;
RAM[16'h6818] = 8'h00;
RAM[16'h6819] = 8'h00;
RAM[16'h681A] = 8'h00;
RAM[16'h681B] = 8'h00;
RAM[16'h681C] = 8'h00;
RAM[16'h681D] = 8'h00;
RAM[16'h681E] = 8'h00;
RAM[16'h681F] = 8'h00;
RAM[16'h6820] = 8'h00;
RAM[16'h6821] = 8'h00;
RAM[16'h6822] = 8'h00;
RAM[16'h6823] = 8'h00;
RAM[16'h6824] = 8'h00;
RAM[16'h6825] = 8'h00;
RAM[16'h6826] = 8'h00;
RAM[16'h6827] = 8'h00;
RAM[16'h6828] = 8'h00;
RAM[16'h6829] = 8'h00;
RAM[16'h682A] = 8'h00;
RAM[16'h682B] = 8'h00;
RAM[16'h682C] = 8'h00;
RAM[16'h682D] = 8'h00;
RAM[16'h682E] = 8'h00;
RAM[16'h682F] = 8'h00;
RAM[16'h6830] = 8'h00;
RAM[16'h6831] = 8'h00;
RAM[16'h6832] = 8'h00;
RAM[16'h6833] = 8'h00;
RAM[16'h6834] = 8'h00;
RAM[16'h6835] = 8'h00;
RAM[16'h6836] = 8'h00;
RAM[16'h6837] = 8'h00;
RAM[16'h6838] = 8'h00;
RAM[16'h6839] = 8'h00;
RAM[16'h683A] = 8'h00;
RAM[16'h683B] = 8'h00;
RAM[16'h683C] = 8'h00;
RAM[16'h683D] = 8'h00;
RAM[16'h683E] = 8'h00;
RAM[16'h683F] = 8'h00;
RAM[16'h6840] = 8'h00;
RAM[16'h6841] = 8'h00;
RAM[16'h6842] = 8'h00;
RAM[16'h6843] = 8'h00;
RAM[16'h6844] = 8'h00;
RAM[16'h6845] = 8'h00;
RAM[16'h6846] = 8'h00;
RAM[16'h6847] = 8'h00;
RAM[16'h6848] = 8'h00;
RAM[16'h6849] = 8'h00;
RAM[16'h684A] = 8'h00;
RAM[16'h684B] = 8'h00;
RAM[16'h684C] = 8'h00;
RAM[16'h684D] = 8'h00;
RAM[16'h684E] = 8'h00;
RAM[16'h684F] = 8'h00;
RAM[16'h6850] = 8'h00;
RAM[16'h6851] = 8'h00;
RAM[16'h6852] = 8'h00;
RAM[16'h6853] = 8'h00;
RAM[16'h6854] = 8'h00;
RAM[16'h6855] = 8'h00;
RAM[16'h6856] = 8'h00;
RAM[16'h6857] = 8'h00;
RAM[16'h6858] = 8'h00;
RAM[16'h6859] = 8'h00;
RAM[16'h685A] = 8'h00;
RAM[16'h685B] = 8'h00;
RAM[16'h685C] = 8'h00;
RAM[16'h685D] = 8'h00;
RAM[16'h685E] = 8'h00;
RAM[16'h685F] = 8'h00;
RAM[16'h6860] = 8'h00;
RAM[16'h6861] = 8'h00;
RAM[16'h6862] = 8'h00;
RAM[16'h6863] = 8'h00;
RAM[16'h6864] = 8'h00;
RAM[16'h6865] = 8'h00;
RAM[16'h6866] = 8'h00;
RAM[16'h6867] = 8'h00;
RAM[16'h6868] = 8'h00;
RAM[16'h6869] = 8'h00;
RAM[16'h686A] = 8'h00;
RAM[16'h686B] = 8'h00;
RAM[16'h686C] = 8'h00;
RAM[16'h686D] = 8'h00;
RAM[16'h686E] = 8'h00;
RAM[16'h686F] = 8'h00;
RAM[16'h6870] = 8'h00;
RAM[16'h6871] = 8'h00;
RAM[16'h6872] = 8'h00;
RAM[16'h6873] = 8'h00;
RAM[16'h6874] = 8'h00;
RAM[16'h6875] = 8'h00;
RAM[16'h6876] = 8'h00;
RAM[16'h6877] = 8'h00;
RAM[16'h6878] = 8'h00;
RAM[16'h6879] = 8'h00;
RAM[16'h687A] = 8'h00;
RAM[16'h687B] = 8'h00;
RAM[16'h687C] = 8'h00;
RAM[16'h687D] = 8'h00;
RAM[16'h687E] = 8'h00;
RAM[16'h687F] = 8'h00;
RAM[16'h6880] = 8'h00;
RAM[16'h6881] = 8'h00;
RAM[16'h6882] = 8'h00;
RAM[16'h6883] = 8'h00;
RAM[16'h6884] = 8'h00;
RAM[16'h6885] = 8'h00;
RAM[16'h6886] = 8'h00;
RAM[16'h6887] = 8'h00;
RAM[16'h6888] = 8'h00;
RAM[16'h6889] = 8'h00;
RAM[16'h688A] = 8'h00;
RAM[16'h688B] = 8'h00;
RAM[16'h688C] = 8'h00;
RAM[16'h688D] = 8'h00;
RAM[16'h688E] = 8'h00;
RAM[16'h688F] = 8'h00;
RAM[16'h6890] = 8'h00;
RAM[16'h6891] = 8'h00;
RAM[16'h6892] = 8'h00;
RAM[16'h6893] = 8'h00;
RAM[16'h6894] = 8'h00;
RAM[16'h6895] = 8'h00;
RAM[16'h6896] = 8'h00;
RAM[16'h6897] = 8'h00;
RAM[16'h6898] = 8'h00;
RAM[16'h6899] = 8'h00;
RAM[16'h689A] = 8'h00;
RAM[16'h689B] = 8'h00;
RAM[16'h689C] = 8'h00;
RAM[16'h689D] = 8'h00;
RAM[16'h689E] = 8'h00;
RAM[16'h689F] = 8'h00;
RAM[16'h68A0] = 8'h00;
RAM[16'h68A1] = 8'h00;
RAM[16'h68A2] = 8'h00;
RAM[16'h68A3] = 8'h00;
RAM[16'h68A4] = 8'h00;
RAM[16'h68A5] = 8'h00;
RAM[16'h68A6] = 8'h00;
RAM[16'h68A7] = 8'h00;
RAM[16'h68A8] = 8'h00;
RAM[16'h68A9] = 8'h00;
RAM[16'h68AA] = 8'h00;
RAM[16'h68AB] = 8'h00;
RAM[16'h68AC] = 8'h00;
RAM[16'h68AD] = 8'h00;
RAM[16'h68AE] = 8'h00;
RAM[16'h68AF] = 8'h00;
RAM[16'h68B0] = 8'h00;
RAM[16'h68B1] = 8'h00;
RAM[16'h68B2] = 8'h00;
RAM[16'h68B3] = 8'h00;
RAM[16'h68B4] = 8'h00;
RAM[16'h68B5] = 8'h00;
RAM[16'h68B6] = 8'h00;
RAM[16'h68B7] = 8'h00;
RAM[16'h68B8] = 8'h00;
RAM[16'h68B9] = 8'h00;
RAM[16'h68BA] = 8'h00;
RAM[16'h68BB] = 8'h00;
RAM[16'h68BC] = 8'h00;
RAM[16'h68BD] = 8'h00;
RAM[16'h68BE] = 8'h00;
RAM[16'h68BF] = 8'h00;
RAM[16'h68C0] = 8'h00;
RAM[16'h68C1] = 8'h00;
RAM[16'h68C2] = 8'h00;
RAM[16'h68C3] = 8'h00;
RAM[16'h68C4] = 8'h00;
RAM[16'h68C5] = 8'h00;
RAM[16'h68C6] = 8'h00;
RAM[16'h68C7] = 8'h00;
RAM[16'h68C8] = 8'h00;
RAM[16'h68C9] = 8'h00;
RAM[16'h68CA] = 8'h00;
RAM[16'h68CB] = 8'h00;
RAM[16'h68CC] = 8'h00;
RAM[16'h68CD] = 8'h00;
RAM[16'h68CE] = 8'h00;
RAM[16'h68CF] = 8'h00;
RAM[16'h68D0] = 8'h00;
RAM[16'h68D1] = 8'h00;
RAM[16'h68D2] = 8'h00;
RAM[16'h68D3] = 8'h00;
RAM[16'h68D4] = 8'h00;
RAM[16'h68D5] = 8'h00;
RAM[16'h68D6] = 8'h00;
RAM[16'h68D7] = 8'h00;
RAM[16'h68D8] = 8'h00;
RAM[16'h68D9] = 8'h00;
RAM[16'h68DA] = 8'h00;
RAM[16'h68DB] = 8'h00;
RAM[16'h68DC] = 8'h00;
RAM[16'h68DD] = 8'h00;
RAM[16'h68DE] = 8'h00;
RAM[16'h68DF] = 8'h00;
RAM[16'h68E0] = 8'h00;
RAM[16'h68E1] = 8'h00;
RAM[16'h68E2] = 8'h00;
RAM[16'h68E3] = 8'h00;
RAM[16'h68E4] = 8'h00;
RAM[16'h68E5] = 8'h00;
RAM[16'h68E6] = 8'h00;
RAM[16'h68E7] = 8'h00;
RAM[16'h68E8] = 8'h00;
RAM[16'h68E9] = 8'h00;
RAM[16'h68EA] = 8'h00;
RAM[16'h68EB] = 8'h00;
RAM[16'h68EC] = 8'h00;
RAM[16'h68ED] = 8'h00;
RAM[16'h68EE] = 8'h00;
RAM[16'h68EF] = 8'h00;
RAM[16'h68F0] = 8'h00;
RAM[16'h68F1] = 8'h00;
RAM[16'h68F2] = 8'h00;
RAM[16'h68F3] = 8'h00;
RAM[16'h68F4] = 8'h00;
RAM[16'h68F5] = 8'h00;
RAM[16'h68F6] = 8'h00;
RAM[16'h68F7] = 8'h00;
RAM[16'h68F8] = 8'h00;
RAM[16'h68F9] = 8'h00;
RAM[16'h68FA] = 8'h00;
RAM[16'h68FB] = 8'h00;
RAM[16'h68FC] = 8'h00;
RAM[16'h68FD] = 8'h00;
RAM[16'h68FE] = 8'h00;
RAM[16'h68FF] = 8'h00;
RAM[16'h6900] = 8'h00;
RAM[16'h6901] = 8'h00;
RAM[16'h6902] = 8'h00;
RAM[16'h6903] = 8'h00;
RAM[16'h6904] = 8'h00;
RAM[16'h6905] = 8'h00;
RAM[16'h6906] = 8'h00;
RAM[16'h6907] = 8'h00;
RAM[16'h6908] = 8'h00;
RAM[16'h6909] = 8'h00;
RAM[16'h690A] = 8'h00;
RAM[16'h690B] = 8'h00;
RAM[16'h690C] = 8'h00;
RAM[16'h690D] = 8'h00;
RAM[16'h690E] = 8'h00;
RAM[16'h690F] = 8'h00;
RAM[16'h6910] = 8'h00;
RAM[16'h6911] = 8'h00;
RAM[16'h6912] = 8'h00;
RAM[16'h6913] = 8'h00;
RAM[16'h6914] = 8'h00;
RAM[16'h6915] = 8'h00;
RAM[16'h6916] = 8'h00;
RAM[16'h6917] = 8'h00;
RAM[16'h6918] = 8'h00;
RAM[16'h6919] = 8'h00;
RAM[16'h691A] = 8'h00;
RAM[16'h691B] = 8'h00;
RAM[16'h691C] = 8'h00;
RAM[16'h691D] = 8'h00;
RAM[16'h691E] = 8'h00;
RAM[16'h691F] = 8'h00;
RAM[16'h6920] = 8'h00;
RAM[16'h6921] = 8'h00;
RAM[16'h6922] = 8'h00;
RAM[16'h6923] = 8'h00;
RAM[16'h6924] = 8'h00;
RAM[16'h6925] = 8'h00;
RAM[16'h6926] = 8'h00;
RAM[16'h6927] = 8'h00;
RAM[16'h6928] = 8'h00;
RAM[16'h6929] = 8'h00;
RAM[16'h692A] = 8'h00;
RAM[16'h692B] = 8'h00;
RAM[16'h692C] = 8'h00;
RAM[16'h692D] = 8'h00;
RAM[16'h692E] = 8'h00;
RAM[16'h692F] = 8'h00;
RAM[16'h6930] = 8'h00;
RAM[16'h6931] = 8'h00;
RAM[16'h6932] = 8'h00;
RAM[16'h6933] = 8'h00;
RAM[16'h6934] = 8'h00;
RAM[16'h6935] = 8'h00;
RAM[16'h6936] = 8'h00;
RAM[16'h6937] = 8'h00;
RAM[16'h6938] = 8'h00;
RAM[16'h6939] = 8'h00;
RAM[16'h693A] = 8'h00;
RAM[16'h693B] = 8'h00;
RAM[16'h693C] = 8'h00;
RAM[16'h693D] = 8'h00;
RAM[16'h693E] = 8'h00;
RAM[16'h693F] = 8'h00;
RAM[16'h6940] = 8'h00;
RAM[16'h6941] = 8'h00;
RAM[16'h6942] = 8'h00;
RAM[16'h6943] = 8'h00;
RAM[16'h6944] = 8'h00;
RAM[16'h6945] = 8'h00;
RAM[16'h6946] = 8'h00;
RAM[16'h6947] = 8'h00;
RAM[16'h6948] = 8'h00;
RAM[16'h6949] = 8'h00;
RAM[16'h694A] = 8'h00;
RAM[16'h694B] = 8'h00;
RAM[16'h694C] = 8'h00;
RAM[16'h694D] = 8'h00;
RAM[16'h694E] = 8'h00;
RAM[16'h694F] = 8'h00;
RAM[16'h6950] = 8'h00;
RAM[16'h6951] = 8'h00;
RAM[16'h6952] = 8'h00;
RAM[16'h6953] = 8'h00;
RAM[16'h6954] = 8'h00;
RAM[16'h6955] = 8'h00;
RAM[16'h6956] = 8'h00;
RAM[16'h6957] = 8'h00;
RAM[16'h6958] = 8'h00;
RAM[16'h6959] = 8'h00;
RAM[16'h695A] = 8'h00;
RAM[16'h695B] = 8'h00;
RAM[16'h695C] = 8'h00;
RAM[16'h695D] = 8'h00;
RAM[16'h695E] = 8'h00;
RAM[16'h695F] = 8'h00;
RAM[16'h6960] = 8'h00;
RAM[16'h6961] = 8'h00;
RAM[16'h6962] = 8'h00;
RAM[16'h6963] = 8'h00;
RAM[16'h6964] = 8'h00;
RAM[16'h6965] = 8'h00;
RAM[16'h6966] = 8'h00;
RAM[16'h6967] = 8'h00;
RAM[16'h6968] = 8'h00;
RAM[16'h6969] = 8'h00;
RAM[16'h696A] = 8'h00;
RAM[16'h696B] = 8'h00;
RAM[16'h696C] = 8'h00;
RAM[16'h696D] = 8'h00;
RAM[16'h696E] = 8'h00;
RAM[16'h696F] = 8'h00;
RAM[16'h6970] = 8'h00;
RAM[16'h6971] = 8'h00;
RAM[16'h6972] = 8'h00;
RAM[16'h6973] = 8'h00;
RAM[16'h6974] = 8'h00;
RAM[16'h6975] = 8'h00;
RAM[16'h6976] = 8'h00;
RAM[16'h6977] = 8'h00;
RAM[16'h6978] = 8'h00;
RAM[16'h6979] = 8'h00;
RAM[16'h697A] = 8'h00;
RAM[16'h697B] = 8'h00;
RAM[16'h697C] = 8'h00;
RAM[16'h697D] = 8'h00;
RAM[16'h697E] = 8'h00;
RAM[16'h697F] = 8'h00;
RAM[16'h6980] = 8'h00;
RAM[16'h6981] = 8'h00;
RAM[16'h6982] = 8'h00;
RAM[16'h6983] = 8'h00;
RAM[16'h6984] = 8'h00;
RAM[16'h6985] = 8'h00;
RAM[16'h6986] = 8'h00;
RAM[16'h6987] = 8'h00;
RAM[16'h6988] = 8'h00;
RAM[16'h6989] = 8'h00;
RAM[16'h698A] = 8'h00;
RAM[16'h698B] = 8'h00;
RAM[16'h698C] = 8'h00;
RAM[16'h698D] = 8'h00;
RAM[16'h698E] = 8'h00;
RAM[16'h698F] = 8'h00;
RAM[16'h6990] = 8'h00;
RAM[16'h6991] = 8'h00;
RAM[16'h6992] = 8'h00;
RAM[16'h6993] = 8'h00;
RAM[16'h6994] = 8'h00;
RAM[16'h6995] = 8'h00;
RAM[16'h6996] = 8'h00;
RAM[16'h6997] = 8'h00;
RAM[16'h6998] = 8'h00;
RAM[16'h6999] = 8'h00;
RAM[16'h699A] = 8'h00;
RAM[16'h699B] = 8'h00;
RAM[16'h699C] = 8'h00;
RAM[16'h699D] = 8'h00;
RAM[16'h699E] = 8'h00;
RAM[16'h699F] = 8'h00;
RAM[16'h69A0] = 8'h00;
RAM[16'h69A1] = 8'h00;
RAM[16'h69A2] = 8'h00;
RAM[16'h69A3] = 8'h00;
RAM[16'h69A4] = 8'h00;
RAM[16'h69A5] = 8'h00;
RAM[16'h69A6] = 8'h00;
RAM[16'h69A7] = 8'h00;
RAM[16'h69A8] = 8'h00;
RAM[16'h69A9] = 8'h00;
RAM[16'h69AA] = 8'h00;
RAM[16'h69AB] = 8'h00;
RAM[16'h69AC] = 8'h00;
RAM[16'h69AD] = 8'h00;
RAM[16'h69AE] = 8'h00;
RAM[16'h69AF] = 8'h00;
RAM[16'h69B0] = 8'h00;
RAM[16'h69B1] = 8'h00;
RAM[16'h69B2] = 8'h00;
RAM[16'h69B3] = 8'h00;
RAM[16'h69B4] = 8'h00;
RAM[16'h69B5] = 8'h00;
RAM[16'h69B6] = 8'h00;
RAM[16'h69B7] = 8'h00;
RAM[16'h69B8] = 8'h00;
RAM[16'h69B9] = 8'h00;
RAM[16'h69BA] = 8'h00;
RAM[16'h69BB] = 8'h00;
RAM[16'h69BC] = 8'h00;
RAM[16'h69BD] = 8'h00;
RAM[16'h69BE] = 8'h00;
RAM[16'h69BF] = 8'h00;
RAM[16'h69C0] = 8'h00;
RAM[16'h69C1] = 8'h00;
RAM[16'h69C2] = 8'h00;
RAM[16'h69C3] = 8'h00;
RAM[16'h69C4] = 8'h00;
RAM[16'h69C5] = 8'h00;
RAM[16'h69C6] = 8'h00;
RAM[16'h69C7] = 8'h00;
RAM[16'h69C8] = 8'h00;
RAM[16'h69C9] = 8'h00;
RAM[16'h69CA] = 8'h00;
RAM[16'h69CB] = 8'h00;
RAM[16'h69CC] = 8'h00;
RAM[16'h69CD] = 8'h00;
RAM[16'h69CE] = 8'h00;
RAM[16'h69CF] = 8'h00;
RAM[16'h69D0] = 8'h00;
RAM[16'h69D1] = 8'h00;
RAM[16'h69D2] = 8'h00;
RAM[16'h69D3] = 8'h00;
RAM[16'h69D4] = 8'h00;
RAM[16'h69D5] = 8'h00;
RAM[16'h69D6] = 8'h00;
RAM[16'h69D7] = 8'h00;
RAM[16'h69D8] = 8'h00;
RAM[16'h69D9] = 8'h00;
RAM[16'h69DA] = 8'h00;
RAM[16'h69DB] = 8'h00;
RAM[16'h69DC] = 8'h00;
RAM[16'h69DD] = 8'h00;
RAM[16'h69DE] = 8'h00;
RAM[16'h69DF] = 8'h00;
RAM[16'h69E0] = 8'h00;
RAM[16'h69E1] = 8'h00;
RAM[16'h69E2] = 8'h00;
RAM[16'h69E3] = 8'h00;
RAM[16'h69E4] = 8'h00;
RAM[16'h69E5] = 8'h00;
RAM[16'h69E6] = 8'h00;
RAM[16'h69E7] = 8'h00;
RAM[16'h69E8] = 8'h00;
RAM[16'h69E9] = 8'h00;
RAM[16'h69EA] = 8'h00;
RAM[16'h69EB] = 8'h00;
RAM[16'h69EC] = 8'h00;
RAM[16'h69ED] = 8'h00;
RAM[16'h69EE] = 8'h00;
RAM[16'h69EF] = 8'h00;
RAM[16'h69F0] = 8'h00;
RAM[16'h69F1] = 8'h00;
RAM[16'h69F2] = 8'h00;
RAM[16'h69F3] = 8'h00;
RAM[16'h69F4] = 8'h00;
RAM[16'h69F5] = 8'h00;
RAM[16'h69F6] = 8'h00;
RAM[16'h69F7] = 8'h00;
RAM[16'h69F8] = 8'h00;
RAM[16'h69F9] = 8'h00;
RAM[16'h69FA] = 8'h00;
RAM[16'h69FB] = 8'h00;
RAM[16'h69FC] = 8'h00;
RAM[16'h69FD] = 8'h00;
RAM[16'h69FE] = 8'h00;
RAM[16'h69FF] = 8'h00;
RAM[16'h6A00] = 8'h00;
RAM[16'h6A01] = 8'h00;
RAM[16'h6A02] = 8'h00;
RAM[16'h6A03] = 8'h00;
RAM[16'h6A04] = 8'h00;
RAM[16'h6A05] = 8'h00;
RAM[16'h6A06] = 8'h00;
RAM[16'h6A07] = 8'h00;
RAM[16'h6A08] = 8'h00;
RAM[16'h6A09] = 8'h00;
RAM[16'h6A0A] = 8'h00;
RAM[16'h6A0B] = 8'h00;
RAM[16'h6A0C] = 8'h00;
RAM[16'h6A0D] = 8'h00;
RAM[16'h6A0E] = 8'h00;
RAM[16'h6A0F] = 8'h00;
RAM[16'h6A10] = 8'h00;
RAM[16'h6A11] = 8'h00;
RAM[16'h6A12] = 8'h00;
RAM[16'h6A13] = 8'h00;
RAM[16'h6A14] = 8'h00;
RAM[16'h6A15] = 8'h00;
RAM[16'h6A16] = 8'h00;
RAM[16'h6A17] = 8'h00;
RAM[16'h6A18] = 8'h00;
RAM[16'h6A19] = 8'h00;
RAM[16'h6A1A] = 8'h00;
RAM[16'h6A1B] = 8'h00;
RAM[16'h6A1C] = 8'h00;
RAM[16'h6A1D] = 8'h00;
RAM[16'h6A1E] = 8'h00;
RAM[16'h6A1F] = 8'h00;
RAM[16'h6A20] = 8'h00;
RAM[16'h6A21] = 8'h00;
RAM[16'h6A22] = 8'h00;
RAM[16'h6A23] = 8'h00;
RAM[16'h6A24] = 8'h00;
RAM[16'h6A25] = 8'h00;
RAM[16'h6A26] = 8'h00;
RAM[16'h6A27] = 8'h00;
RAM[16'h6A28] = 8'h00;
RAM[16'h6A29] = 8'h00;
RAM[16'h6A2A] = 8'h00;
RAM[16'h6A2B] = 8'h00;
RAM[16'h6A2C] = 8'h00;
RAM[16'h6A2D] = 8'h00;
RAM[16'h6A2E] = 8'h00;
RAM[16'h6A2F] = 8'h00;
RAM[16'h6A30] = 8'h00;
RAM[16'h6A31] = 8'h00;
RAM[16'h6A32] = 8'h00;
RAM[16'h6A33] = 8'h00;
RAM[16'h6A34] = 8'h00;
RAM[16'h6A35] = 8'h00;
RAM[16'h6A36] = 8'h00;
RAM[16'h6A37] = 8'h00;
RAM[16'h6A38] = 8'h00;
RAM[16'h6A39] = 8'h00;
RAM[16'h6A3A] = 8'h00;
RAM[16'h6A3B] = 8'h00;
RAM[16'h6A3C] = 8'h00;
RAM[16'h6A3D] = 8'h00;
RAM[16'h6A3E] = 8'h00;
RAM[16'h6A3F] = 8'h00;
RAM[16'h6A40] = 8'h00;
RAM[16'h6A41] = 8'h00;
RAM[16'h6A42] = 8'h00;
RAM[16'h6A43] = 8'h00;
RAM[16'h6A44] = 8'h00;
RAM[16'h6A45] = 8'h00;
RAM[16'h6A46] = 8'h00;
RAM[16'h6A47] = 8'h00;
RAM[16'h6A48] = 8'h00;
RAM[16'h6A49] = 8'h00;
RAM[16'h6A4A] = 8'h00;
RAM[16'h6A4B] = 8'h00;
RAM[16'h6A4C] = 8'h00;
RAM[16'h6A4D] = 8'h00;
RAM[16'h6A4E] = 8'h00;
RAM[16'h6A4F] = 8'h00;
RAM[16'h6A50] = 8'h00;
RAM[16'h6A51] = 8'h00;
RAM[16'h6A52] = 8'h00;
RAM[16'h6A53] = 8'h00;
RAM[16'h6A54] = 8'h00;
RAM[16'h6A55] = 8'h00;
RAM[16'h6A56] = 8'h00;
RAM[16'h6A57] = 8'h00;
RAM[16'h6A58] = 8'h00;
RAM[16'h6A59] = 8'h00;
RAM[16'h6A5A] = 8'h00;
RAM[16'h6A5B] = 8'h00;
RAM[16'h6A5C] = 8'h00;
RAM[16'h6A5D] = 8'h00;
RAM[16'h6A5E] = 8'h00;
RAM[16'h6A5F] = 8'h00;
RAM[16'h6A60] = 8'h00;
RAM[16'h6A61] = 8'h00;
RAM[16'h6A62] = 8'h00;
RAM[16'h6A63] = 8'h00;
RAM[16'h6A64] = 8'h00;
RAM[16'h6A65] = 8'h00;
RAM[16'h6A66] = 8'h00;
RAM[16'h6A67] = 8'h00;
RAM[16'h6A68] = 8'h00;
RAM[16'h6A69] = 8'h00;
RAM[16'h6A6A] = 8'h00;
RAM[16'h6A6B] = 8'h00;
RAM[16'h6A6C] = 8'h00;
RAM[16'h6A6D] = 8'h00;
RAM[16'h6A6E] = 8'h00;
RAM[16'h6A6F] = 8'h00;
RAM[16'h6A70] = 8'h00;
RAM[16'h6A71] = 8'h00;
RAM[16'h6A72] = 8'h00;
RAM[16'h6A73] = 8'h00;
RAM[16'h6A74] = 8'h00;
RAM[16'h6A75] = 8'h00;
RAM[16'h6A76] = 8'h00;
RAM[16'h6A77] = 8'h00;
RAM[16'h6A78] = 8'h00;
RAM[16'h6A79] = 8'h00;
RAM[16'h6A7A] = 8'h00;
RAM[16'h6A7B] = 8'h00;
RAM[16'h6A7C] = 8'h00;
RAM[16'h6A7D] = 8'h00;
RAM[16'h6A7E] = 8'h00;
RAM[16'h6A7F] = 8'h00;
RAM[16'h6A80] = 8'h00;
RAM[16'h6A81] = 8'h00;
RAM[16'h6A82] = 8'h00;
RAM[16'h6A83] = 8'h00;
RAM[16'h6A84] = 8'h00;
RAM[16'h6A85] = 8'h00;
RAM[16'h6A86] = 8'h00;
RAM[16'h6A87] = 8'h00;
RAM[16'h6A88] = 8'h00;
RAM[16'h6A89] = 8'h00;
RAM[16'h6A8A] = 8'h00;
RAM[16'h6A8B] = 8'h00;
RAM[16'h6A8C] = 8'h00;
RAM[16'h6A8D] = 8'h00;
RAM[16'h6A8E] = 8'h00;
RAM[16'h6A8F] = 8'h00;
RAM[16'h6A90] = 8'h00;
RAM[16'h6A91] = 8'h00;
RAM[16'h6A92] = 8'h00;
RAM[16'h6A93] = 8'h00;
RAM[16'h6A94] = 8'h00;
RAM[16'h6A95] = 8'h00;
RAM[16'h6A96] = 8'h00;
RAM[16'h6A97] = 8'h00;
RAM[16'h6A98] = 8'h00;
RAM[16'h6A99] = 8'h00;
RAM[16'h6A9A] = 8'h00;
RAM[16'h6A9B] = 8'h00;
RAM[16'h6A9C] = 8'h00;
RAM[16'h6A9D] = 8'h00;
RAM[16'h6A9E] = 8'h00;
RAM[16'h6A9F] = 8'h00;
RAM[16'h6AA0] = 8'h00;
RAM[16'h6AA1] = 8'h00;
RAM[16'h6AA2] = 8'h00;
RAM[16'h6AA3] = 8'h00;
RAM[16'h6AA4] = 8'h00;
RAM[16'h6AA5] = 8'h00;
RAM[16'h6AA6] = 8'h00;
RAM[16'h6AA7] = 8'h00;
RAM[16'h6AA8] = 8'h00;
RAM[16'h6AA9] = 8'h00;
RAM[16'h6AAA] = 8'h00;
RAM[16'h6AAB] = 8'h00;
RAM[16'h6AAC] = 8'h00;
RAM[16'h6AAD] = 8'h00;
RAM[16'h6AAE] = 8'h00;
RAM[16'h6AAF] = 8'h00;
RAM[16'h6AB0] = 8'h00;
RAM[16'h6AB1] = 8'h00;
RAM[16'h6AB2] = 8'h00;
RAM[16'h6AB3] = 8'h00;
RAM[16'h6AB4] = 8'h00;
RAM[16'h6AB5] = 8'h00;
RAM[16'h6AB6] = 8'h00;
RAM[16'h6AB7] = 8'h00;
RAM[16'h6AB8] = 8'h00;
RAM[16'h6AB9] = 8'h00;
RAM[16'h6ABA] = 8'h00;
RAM[16'h6ABB] = 8'h00;
RAM[16'h6ABC] = 8'h00;
RAM[16'h6ABD] = 8'h00;
RAM[16'h6ABE] = 8'h00;
RAM[16'h6ABF] = 8'h00;
RAM[16'h6AC0] = 8'h00;
RAM[16'h6AC1] = 8'h00;
RAM[16'h6AC2] = 8'h00;
RAM[16'h6AC3] = 8'h00;
RAM[16'h6AC4] = 8'h00;
RAM[16'h6AC5] = 8'h00;
RAM[16'h6AC6] = 8'h00;
RAM[16'h6AC7] = 8'h00;
RAM[16'h6AC8] = 8'h00;
RAM[16'h6AC9] = 8'h00;
RAM[16'h6ACA] = 8'h00;
RAM[16'h6ACB] = 8'h00;
RAM[16'h6ACC] = 8'h00;
RAM[16'h6ACD] = 8'h00;
RAM[16'h6ACE] = 8'h00;
RAM[16'h6ACF] = 8'h00;
RAM[16'h6AD0] = 8'h00;
RAM[16'h6AD1] = 8'h00;
RAM[16'h6AD2] = 8'h00;
RAM[16'h6AD3] = 8'h00;
RAM[16'h6AD4] = 8'h00;
RAM[16'h6AD5] = 8'h00;
RAM[16'h6AD6] = 8'h00;
RAM[16'h6AD7] = 8'h00;
RAM[16'h6AD8] = 8'h00;
RAM[16'h6AD9] = 8'h00;
RAM[16'h6ADA] = 8'h00;
RAM[16'h6ADB] = 8'h00;
RAM[16'h6ADC] = 8'h00;
RAM[16'h6ADD] = 8'h00;
RAM[16'h6ADE] = 8'h00;
RAM[16'h6ADF] = 8'h00;
RAM[16'h6AE0] = 8'h00;
RAM[16'h6AE1] = 8'h00;
RAM[16'h6AE2] = 8'h00;
RAM[16'h6AE3] = 8'h00;
RAM[16'h6AE4] = 8'h00;
RAM[16'h6AE5] = 8'h00;
RAM[16'h6AE6] = 8'h00;
RAM[16'h6AE7] = 8'h00;
RAM[16'h6AE8] = 8'h00;
RAM[16'h6AE9] = 8'h00;
RAM[16'h6AEA] = 8'h00;
RAM[16'h6AEB] = 8'h00;
RAM[16'h6AEC] = 8'h00;
RAM[16'h6AED] = 8'h00;
RAM[16'h6AEE] = 8'h00;
RAM[16'h6AEF] = 8'h00;
RAM[16'h6AF0] = 8'h00;
RAM[16'h6AF1] = 8'h00;
RAM[16'h6AF2] = 8'h00;
RAM[16'h6AF3] = 8'h00;
RAM[16'h6AF4] = 8'h00;
RAM[16'h6AF5] = 8'h00;
RAM[16'h6AF6] = 8'h00;
RAM[16'h6AF7] = 8'h00;
RAM[16'h6AF8] = 8'h00;
RAM[16'h6AF9] = 8'h00;
RAM[16'h6AFA] = 8'h00;
RAM[16'h6AFB] = 8'h00;
RAM[16'h6AFC] = 8'h00;
RAM[16'h6AFD] = 8'h00;
RAM[16'h6AFE] = 8'h00;
RAM[16'h6AFF] = 8'h00;
RAM[16'h6B00] = 8'h00;
RAM[16'h6B01] = 8'h00;
RAM[16'h6B02] = 8'h00;
RAM[16'h6B03] = 8'h00;
RAM[16'h6B04] = 8'h00;
RAM[16'h6B05] = 8'h00;
RAM[16'h6B06] = 8'h00;
RAM[16'h6B07] = 8'h00;
RAM[16'h6B08] = 8'h00;
RAM[16'h6B09] = 8'h00;
RAM[16'h6B0A] = 8'h00;
RAM[16'h6B0B] = 8'h00;
RAM[16'h6B0C] = 8'h00;
RAM[16'h6B0D] = 8'h00;
RAM[16'h6B0E] = 8'h00;
RAM[16'h6B0F] = 8'h00;
RAM[16'h6B10] = 8'h00;
RAM[16'h6B11] = 8'h00;
RAM[16'h6B12] = 8'h00;
RAM[16'h6B13] = 8'h00;
RAM[16'h6B14] = 8'h00;
RAM[16'h6B15] = 8'h00;
RAM[16'h6B16] = 8'h00;
RAM[16'h6B17] = 8'h00;
RAM[16'h6B18] = 8'h00;
RAM[16'h6B19] = 8'h00;
RAM[16'h6B1A] = 8'h00;
RAM[16'h6B1B] = 8'h00;
RAM[16'h6B1C] = 8'h00;
RAM[16'h6B1D] = 8'h00;
RAM[16'h6B1E] = 8'h00;
RAM[16'h6B1F] = 8'h00;
RAM[16'h6B20] = 8'h00;
RAM[16'h6B21] = 8'h00;
RAM[16'h6B22] = 8'h00;
RAM[16'h6B23] = 8'h00;
RAM[16'h6B24] = 8'h00;
RAM[16'h6B25] = 8'h00;
RAM[16'h6B26] = 8'h00;
RAM[16'h6B27] = 8'h00;
RAM[16'h6B28] = 8'h00;
RAM[16'h6B29] = 8'h00;
RAM[16'h6B2A] = 8'h00;
RAM[16'h6B2B] = 8'h00;
RAM[16'h6B2C] = 8'h00;
RAM[16'h6B2D] = 8'h00;
RAM[16'h6B2E] = 8'h00;
RAM[16'h6B2F] = 8'h00;
RAM[16'h6B30] = 8'h00;
RAM[16'h6B31] = 8'h00;
RAM[16'h6B32] = 8'h00;
RAM[16'h6B33] = 8'h00;
RAM[16'h6B34] = 8'h00;
RAM[16'h6B35] = 8'h00;
RAM[16'h6B36] = 8'h00;
RAM[16'h6B37] = 8'h00;
RAM[16'h6B38] = 8'h00;
RAM[16'h6B39] = 8'h00;
RAM[16'h6B3A] = 8'h00;
RAM[16'h6B3B] = 8'h00;
RAM[16'h6B3C] = 8'h00;
RAM[16'h6B3D] = 8'h00;
RAM[16'h6B3E] = 8'h00;
RAM[16'h6B3F] = 8'h00;
RAM[16'h6B40] = 8'h00;
RAM[16'h6B41] = 8'h00;
RAM[16'h6B42] = 8'h00;
RAM[16'h6B43] = 8'h00;
RAM[16'h6B44] = 8'h00;
RAM[16'h6B45] = 8'h00;
RAM[16'h6B46] = 8'h00;
RAM[16'h6B47] = 8'h00;
RAM[16'h6B48] = 8'h00;
RAM[16'h6B49] = 8'h00;
RAM[16'h6B4A] = 8'h00;
RAM[16'h6B4B] = 8'h00;
RAM[16'h6B4C] = 8'h00;
RAM[16'h6B4D] = 8'h00;
RAM[16'h6B4E] = 8'h00;
RAM[16'h6B4F] = 8'h00;
RAM[16'h6B50] = 8'h00;
RAM[16'h6B51] = 8'h00;
RAM[16'h6B52] = 8'h00;
RAM[16'h6B53] = 8'h00;
RAM[16'h6B54] = 8'h00;
RAM[16'h6B55] = 8'h00;
RAM[16'h6B56] = 8'h00;
RAM[16'h6B57] = 8'h00;
RAM[16'h6B58] = 8'h00;
RAM[16'h6B59] = 8'h00;
RAM[16'h6B5A] = 8'h00;
RAM[16'h6B5B] = 8'h00;
RAM[16'h6B5C] = 8'h00;
RAM[16'h6B5D] = 8'h00;
RAM[16'h6B5E] = 8'h00;
RAM[16'h6B5F] = 8'h00;
RAM[16'h6B60] = 8'h00;
RAM[16'h6B61] = 8'h00;
RAM[16'h6B62] = 8'h00;
RAM[16'h6B63] = 8'h00;
RAM[16'h6B64] = 8'h00;
RAM[16'h6B65] = 8'h00;
RAM[16'h6B66] = 8'h00;
RAM[16'h6B67] = 8'h00;
RAM[16'h6B68] = 8'h00;
RAM[16'h6B69] = 8'h00;
RAM[16'h6B6A] = 8'h00;
RAM[16'h6B6B] = 8'h00;
RAM[16'h6B6C] = 8'h00;
RAM[16'h6B6D] = 8'h00;
RAM[16'h6B6E] = 8'h00;
RAM[16'h6B6F] = 8'h00;
RAM[16'h6B70] = 8'h00;
RAM[16'h6B71] = 8'h00;
RAM[16'h6B72] = 8'h00;
RAM[16'h6B73] = 8'h00;
RAM[16'h6B74] = 8'h00;
RAM[16'h6B75] = 8'h00;
RAM[16'h6B76] = 8'h00;
RAM[16'h6B77] = 8'h00;
RAM[16'h6B78] = 8'h00;
RAM[16'h6B79] = 8'h00;
RAM[16'h6B7A] = 8'h00;
RAM[16'h6B7B] = 8'h00;
RAM[16'h6B7C] = 8'h00;
RAM[16'h6B7D] = 8'h00;
RAM[16'h6B7E] = 8'h00;
RAM[16'h6B7F] = 8'h00;
RAM[16'h6B80] = 8'h00;
RAM[16'h6B81] = 8'h00;
RAM[16'h6B82] = 8'h00;
RAM[16'h6B83] = 8'h00;
RAM[16'h6B84] = 8'h00;
RAM[16'h6B85] = 8'h00;
RAM[16'h6B86] = 8'h00;
RAM[16'h6B87] = 8'h00;
RAM[16'h6B88] = 8'h00;
RAM[16'h6B89] = 8'h00;
RAM[16'h6B8A] = 8'h00;
RAM[16'h6B8B] = 8'h00;
RAM[16'h6B8C] = 8'h00;
RAM[16'h6B8D] = 8'h00;
RAM[16'h6B8E] = 8'h00;
RAM[16'h6B8F] = 8'h00;
RAM[16'h6B90] = 8'h00;
RAM[16'h6B91] = 8'h00;
RAM[16'h6B92] = 8'h00;
RAM[16'h6B93] = 8'h00;
RAM[16'h6B94] = 8'h00;
RAM[16'h6B95] = 8'h00;
RAM[16'h6B96] = 8'h00;
RAM[16'h6B97] = 8'h00;
RAM[16'h6B98] = 8'h00;
RAM[16'h6B99] = 8'h00;
RAM[16'h6B9A] = 8'h00;
RAM[16'h6B9B] = 8'h00;
RAM[16'h6B9C] = 8'h00;
RAM[16'h6B9D] = 8'h00;
RAM[16'h6B9E] = 8'h00;
RAM[16'h6B9F] = 8'h00;
RAM[16'h6BA0] = 8'h00;
RAM[16'h6BA1] = 8'h00;
RAM[16'h6BA2] = 8'h00;
RAM[16'h6BA3] = 8'h00;
RAM[16'h6BA4] = 8'h00;
RAM[16'h6BA5] = 8'h00;
RAM[16'h6BA6] = 8'h00;
RAM[16'h6BA7] = 8'h00;
RAM[16'h6BA8] = 8'h00;
RAM[16'h6BA9] = 8'h00;
RAM[16'h6BAA] = 8'h00;
RAM[16'h6BAB] = 8'h00;
RAM[16'h6BAC] = 8'h00;
RAM[16'h6BAD] = 8'h00;
RAM[16'h6BAE] = 8'h00;
RAM[16'h6BAF] = 8'h00;
RAM[16'h6BB0] = 8'h00;
RAM[16'h6BB1] = 8'h00;
RAM[16'h6BB2] = 8'h00;
RAM[16'h6BB3] = 8'h00;
RAM[16'h6BB4] = 8'h00;
RAM[16'h6BB5] = 8'h00;
RAM[16'h6BB6] = 8'h00;
RAM[16'h6BB7] = 8'h00;
RAM[16'h6BB8] = 8'h00;
RAM[16'h6BB9] = 8'h00;
RAM[16'h6BBA] = 8'h00;
RAM[16'h6BBB] = 8'h00;
RAM[16'h6BBC] = 8'h00;
RAM[16'h6BBD] = 8'h00;
RAM[16'h6BBE] = 8'h00;
RAM[16'h6BBF] = 8'h00;
RAM[16'h6BC0] = 8'h00;
RAM[16'h6BC1] = 8'h00;
RAM[16'h6BC2] = 8'h00;
RAM[16'h6BC3] = 8'h00;
RAM[16'h6BC4] = 8'h00;
RAM[16'h6BC5] = 8'h00;
RAM[16'h6BC6] = 8'h00;
RAM[16'h6BC7] = 8'h00;
RAM[16'h6BC8] = 8'h00;
RAM[16'h6BC9] = 8'h00;
RAM[16'h6BCA] = 8'h00;
RAM[16'h6BCB] = 8'h00;
RAM[16'h6BCC] = 8'h00;
RAM[16'h6BCD] = 8'h00;
RAM[16'h6BCE] = 8'h00;
RAM[16'h6BCF] = 8'h00;
RAM[16'h6BD0] = 8'h00;
RAM[16'h6BD1] = 8'h00;
RAM[16'h6BD2] = 8'h00;
RAM[16'h6BD3] = 8'h00;
RAM[16'h6BD4] = 8'h00;
RAM[16'h6BD5] = 8'h00;
RAM[16'h6BD6] = 8'h00;
RAM[16'h6BD7] = 8'h00;
RAM[16'h6BD8] = 8'h00;
RAM[16'h6BD9] = 8'h00;
RAM[16'h6BDA] = 8'h00;
RAM[16'h6BDB] = 8'h00;
RAM[16'h6BDC] = 8'h00;
RAM[16'h6BDD] = 8'h00;
RAM[16'h6BDE] = 8'h00;
RAM[16'h6BDF] = 8'h00;
RAM[16'h6BE0] = 8'h00;
RAM[16'h6BE1] = 8'h00;
RAM[16'h6BE2] = 8'h00;
RAM[16'h6BE3] = 8'h00;
RAM[16'h6BE4] = 8'h00;
RAM[16'h6BE5] = 8'h00;
RAM[16'h6BE6] = 8'h00;
RAM[16'h6BE7] = 8'h00;
RAM[16'h6BE8] = 8'h00;
RAM[16'h6BE9] = 8'h00;
RAM[16'h6BEA] = 8'h00;
RAM[16'h6BEB] = 8'h00;
RAM[16'h6BEC] = 8'h00;
RAM[16'h6BED] = 8'h00;
RAM[16'h6BEE] = 8'h00;
RAM[16'h6BEF] = 8'h00;
RAM[16'h6BF0] = 8'h00;
RAM[16'h6BF1] = 8'h00;
RAM[16'h6BF2] = 8'h00;
RAM[16'h6BF3] = 8'h00;
RAM[16'h6BF4] = 8'h00;
RAM[16'h6BF5] = 8'h00;
RAM[16'h6BF6] = 8'h00;
RAM[16'h6BF7] = 8'h00;
RAM[16'h6BF8] = 8'h00;
RAM[16'h6BF9] = 8'h00;
RAM[16'h6BFA] = 8'h00;
RAM[16'h6BFB] = 8'h00;
RAM[16'h6BFC] = 8'h00;
RAM[16'h6BFD] = 8'h00;
RAM[16'h6BFE] = 8'h00;
RAM[16'h6BFF] = 8'h00;
RAM[16'h6C00] = 8'h00;
RAM[16'h6C01] = 8'h00;
RAM[16'h6C02] = 8'h00;
RAM[16'h6C03] = 8'h00;
RAM[16'h6C04] = 8'h00;
RAM[16'h6C05] = 8'h00;
RAM[16'h6C06] = 8'h00;
RAM[16'h6C07] = 8'h00;
RAM[16'h6C08] = 8'h00;
RAM[16'h6C09] = 8'h00;
RAM[16'h6C0A] = 8'h00;
RAM[16'h6C0B] = 8'h00;
RAM[16'h6C0C] = 8'h00;
RAM[16'h6C0D] = 8'h00;
RAM[16'h6C0E] = 8'h00;
RAM[16'h6C0F] = 8'h00;
RAM[16'h6C10] = 8'h00;
RAM[16'h6C11] = 8'h00;
RAM[16'h6C12] = 8'h00;
RAM[16'h6C13] = 8'h00;
RAM[16'h6C14] = 8'h00;
RAM[16'h6C15] = 8'h00;
RAM[16'h6C16] = 8'h00;
RAM[16'h6C17] = 8'h00;
RAM[16'h6C18] = 8'h00;
RAM[16'h6C19] = 8'h00;
RAM[16'h6C1A] = 8'h00;
RAM[16'h6C1B] = 8'h00;
RAM[16'h6C1C] = 8'h00;
RAM[16'h6C1D] = 8'h00;
RAM[16'h6C1E] = 8'h00;
RAM[16'h6C1F] = 8'h00;
RAM[16'h6C20] = 8'h00;
RAM[16'h6C21] = 8'h00;
RAM[16'h6C22] = 8'h00;
RAM[16'h6C23] = 8'h00;
RAM[16'h6C24] = 8'h00;
RAM[16'h6C25] = 8'h00;
RAM[16'h6C26] = 8'h00;
RAM[16'h6C27] = 8'h00;
RAM[16'h6C28] = 8'h00;
RAM[16'h6C29] = 8'h00;
RAM[16'h6C2A] = 8'h00;
RAM[16'h6C2B] = 8'h00;
RAM[16'h6C2C] = 8'h00;
RAM[16'h6C2D] = 8'h00;
RAM[16'h6C2E] = 8'h00;
RAM[16'h6C2F] = 8'h00;
RAM[16'h6C30] = 8'h00;
RAM[16'h6C31] = 8'h00;
RAM[16'h6C32] = 8'h00;
RAM[16'h6C33] = 8'h00;
RAM[16'h6C34] = 8'h00;
RAM[16'h6C35] = 8'h00;
RAM[16'h6C36] = 8'h00;
RAM[16'h6C37] = 8'h00;
RAM[16'h6C38] = 8'h00;
RAM[16'h6C39] = 8'h00;
RAM[16'h6C3A] = 8'h00;
RAM[16'h6C3B] = 8'h00;
RAM[16'h6C3C] = 8'h00;
RAM[16'h6C3D] = 8'h00;
RAM[16'h6C3E] = 8'h00;
RAM[16'h6C3F] = 8'h00;
RAM[16'h6C40] = 8'h00;
RAM[16'h6C41] = 8'h00;
RAM[16'h6C42] = 8'h00;
RAM[16'h6C43] = 8'h00;
RAM[16'h6C44] = 8'h00;
RAM[16'h6C45] = 8'h00;
RAM[16'h6C46] = 8'h00;
RAM[16'h6C47] = 8'h00;
RAM[16'h6C48] = 8'h00;
RAM[16'h6C49] = 8'h00;
RAM[16'h6C4A] = 8'h00;
RAM[16'h6C4B] = 8'h00;
RAM[16'h6C4C] = 8'h00;
RAM[16'h6C4D] = 8'h00;
RAM[16'h6C4E] = 8'h00;
RAM[16'h6C4F] = 8'h00;
RAM[16'h6C50] = 8'h00;
RAM[16'h6C51] = 8'h00;
RAM[16'h6C52] = 8'h00;
RAM[16'h6C53] = 8'h00;
RAM[16'h6C54] = 8'h00;
RAM[16'h6C55] = 8'h00;
RAM[16'h6C56] = 8'h00;
RAM[16'h6C57] = 8'h00;
RAM[16'h6C58] = 8'h00;
RAM[16'h6C59] = 8'h00;
RAM[16'h6C5A] = 8'h00;
RAM[16'h6C5B] = 8'h00;
RAM[16'h6C5C] = 8'h00;
RAM[16'h6C5D] = 8'h00;
RAM[16'h6C5E] = 8'h00;
RAM[16'h6C5F] = 8'h00;
RAM[16'h6C60] = 8'h00;
RAM[16'h6C61] = 8'h00;
RAM[16'h6C62] = 8'h00;
RAM[16'h6C63] = 8'h00;
RAM[16'h6C64] = 8'h00;
RAM[16'h6C65] = 8'h00;
RAM[16'h6C66] = 8'h00;
RAM[16'h6C67] = 8'h00;
RAM[16'h6C68] = 8'h00;
RAM[16'h6C69] = 8'h00;
RAM[16'h6C6A] = 8'h00;
RAM[16'h6C6B] = 8'h00;
RAM[16'h6C6C] = 8'h00;
RAM[16'h6C6D] = 8'h00;
RAM[16'h6C6E] = 8'h00;
RAM[16'h6C6F] = 8'h00;
RAM[16'h6C70] = 8'h00;
RAM[16'h6C71] = 8'h00;
RAM[16'h6C72] = 8'h00;
RAM[16'h6C73] = 8'h00;
RAM[16'h6C74] = 8'h00;
RAM[16'h6C75] = 8'h00;
RAM[16'h6C76] = 8'h00;
RAM[16'h6C77] = 8'h00;
RAM[16'h6C78] = 8'h00;
RAM[16'h6C79] = 8'h00;
RAM[16'h6C7A] = 8'h00;
RAM[16'h6C7B] = 8'h00;
RAM[16'h6C7C] = 8'h00;
RAM[16'h6C7D] = 8'h00;
RAM[16'h6C7E] = 8'h00;
RAM[16'h6C7F] = 8'h00;
RAM[16'h6C80] = 8'h00;
RAM[16'h6C81] = 8'h00;
RAM[16'h6C82] = 8'h00;
RAM[16'h6C83] = 8'h00;
RAM[16'h6C84] = 8'h00;
RAM[16'h6C85] = 8'h00;
RAM[16'h6C86] = 8'h00;
RAM[16'h6C87] = 8'h00;
RAM[16'h6C88] = 8'h00;
RAM[16'h6C89] = 8'h00;
RAM[16'h6C8A] = 8'h00;
RAM[16'h6C8B] = 8'h00;
RAM[16'h6C8C] = 8'h00;
RAM[16'h6C8D] = 8'h00;
RAM[16'h6C8E] = 8'h00;
RAM[16'h6C8F] = 8'h00;
RAM[16'h6C90] = 8'h00;
RAM[16'h6C91] = 8'h00;
RAM[16'h6C92] = 8'h00;
RAM[16'h6C93] = 8'h00;
RAM[16'h6C94] = 8'h00;
RAM[16'h6C95] = 8'h00;
RAM[16'h6C96] = 8'h00;
RAM[16'h6C97] = 8'h00;
RAM[16'h6C98] = 8'h00;
RAM[16'h6C99] = 8'h00;
RAM[16'h6C9A] = 8'h00;
RAM[16'h6C9B] = 8'h00;
RAM[16'h6C9C] = 8'h00;
RAM[16'h6C9D] = 8'h00;
RAM[16'h6C9E] = 8'h00;
RAM[16'h6C9F] = 8'h00;
RAM[16'h6CA0] = 8'h00;
RAM[16'h6CA1] = 8'h00;
RAM[16'h6CA2] = 8'h00;
RAM[16'h6CA3] = 8'h00;
RAM[16'h6CA4] = 8'h00;
RAM[16'h6CA5] = 8'h00;
RAM[16'h6CA6] = 8'h00;
RAM[16'h6CA7] = 8'h00;
RAM[16'h6CA8] = 8'h00;
RAM[16'h6CA9] = 8'h00;
RAM[16'h6CAA] = 8'h00;
RAM[16'h6CAB] = 8'h00;
RAM[16'h6CAC] = 8'h00;
RAM[16'h6CAD] = 8'h00;
RAM[16'h6CAE] = 8'h00;
RAM[16'h6CAF] = 8'h00;
RAM[16'h6CB0] = 8'h00;
RAM[16'h6CB1] = 8'h00;
RAM[16'h6CB2] = 8'h00;
RAM[16'h6CB3] = 8'h00;
RAM[16'h6CB4] = 8'h00;
RAM[16'h6CB5] = 8'h00;
RAM[16'h6CB6] = 8'h00;
RAM[16'h6CB7] = 8'h00;
RAM[16'h6CB8] = 8'h00;
RAM[16'h6CB9] = 8'h00;
RAM[16'h6CBA] = 8'h00;
RAM[16'h6CBB] = 8'h00;
RAM[16'h6CBC] = 8'h00;
RAM[16'h6CBD] = 8'h00;
RAM[16'h6CBE] = 8'h00;
RAM[16'h6CBF] = 8'h00;
RAM[16'h6CC0] = 8'h00;
RAM[16'h6CC1] = 8'h00;
RAM[16'h6CC2] = 8'h00;
RAM[16'h6CC3] = 8'h00;
RAM[16'h6CC4] = 8'h00;
RAM[16'h6CC5] = 8'h00;
RAM[16'h6CC6] = 8'h00;
RAM[16'h6CC7] = 8'h00;
RAM[16'h6CC8] = 8'h00;
RAM[16'h6CC9] = 8'h00;
RAM[16'h6CCA] = 8'h00;
RAM[16'h6CCB] = 8'h00;
RAM[16'h6CCC] = 8'h00;
RAM[16'h6CCD] = 8'h00;
RAM[16'h6CCE] = 8'h00;
RAM[16'h6CCF] = 8'h00;
RAM[16'h6CD0] = 8'h00;
RAM[16'h6CD1] = 8'h00;
RAM[16'h6CD2] = 8'h00;
RAM[16'h6CD3] = 8'h00;
RAM[16'h6CD4] = 8'h00;
RAM[16'h6CD5] = 8'h00;
RAM[16'h6CD6] = 8'h00;
RAM[16'h6CD7] = 8'h00;
RAM[16'h6CD8] = 8'h00;
RAM[16'h6CD9] = 8'h00;
RAM[16'h6CDA] = 8'h00;
RAM[16'h6CDB] = 8'h00;
RAM[16'h6CDC] = 8'h00;
RAM[16'h6CDD] = 8'h00;
RAM[16'h6CDE] = 8'h00;
RAM[16'h6CDF] = 8'h00;
RAM[16'h6CE0] = 8'h00;
RAM[16'h6CE1] = 8'h00;
RAM[16'h6CE2] = 8'h00;
RAM[16'h6CE3] = 8'h00;
RAM[16'h6CE4] = 8'h00;
RAM[16'h6CE5] = 8'h00;
RAM[16'h6CE6] = 8'h00;
RAM[16'h6CE7] = 8'h00;
RAM[16'h6CE8] = 8'h00;
RAM[16'h6CE9] = 8'h00;
RAM[16'h6CEA] = 8'h00;
RAM[16'h6CEB] = 8'h00;
RAM[16'h6CEC] = 8'h00;
RAM[16'h6CED] = 8'h00;
RAM[16'h6CEE] = 8'h00;
RAM[16'h6CEF] = 8'h00;
RAM[16'h6CF0] = 8'h00;
RAM[16'h6CF1] = 8'h00;
RAM[16'h6CF2] = 8'h00;
RAM[16'h6CF3] = 8'h00;
RAM[16'h6CF4] = 8'h00;
RAM[16'h6CF5] = 8'h00;
RAM[16'h6CF6] = 8'h00;
RAM[16'h6CF7] = 8'h00;
RAM[16'h6CF8] = 8'h00;
RAM[16'h6CF9] = 8'h00;
RAM[16'h6CFA] = 8'h00;
RAM[16'h6CFB] = 8'h00;
RAM[16'h6CFC] = 8'h00;
RAM[16'h6CFD] = 8'h00;
RAM[16'h6CFE] = 8'h00;
RAM[16'h6CFF] = 8'h00;
RAM[16'h6D00] = 8'h00;
RAM[16'h6D01] = 8'h00;
RAM[16'h6D02] = 8'h00;
RAM[16'h6D03] = 8'h00;
RAM[16'h6D04] = 8'h00;
RAM[16'h6D05] = 8'h00;
RAM[16'h6D06] = 8'h00;
RAM[16'h6D07] = 8'h00;
RAM[16'h6D08] = 8'h00;
RAM[16'h6D09] = 8'h00;
RAM[16'h6D0A] = 8'h00;
RAM[16'h6D0B] = 8'h00;
RAM[16'h6D0C] = 8'h00;
RAM[16'h6D0D] = 8'h00;
RAM[16'h6D0E] = 8'h00;
RAM[16'h6D0F] = 8'h00;
RAM[16'h6D10] = 8'h00;
RAM[16'h6D11] = 8'h00;
RAM[16'h6D12] = 8'h00;
RAM[16'h6D13] = 8'h00;
RAM[16'h6D14] = 8'h00;
RAM[16'h6D15] = 8'h00;
RAM[16'h6D16] = 8'h00;
RAM[16'h6D17] = 8'h00;
RAM[16'h6D18] = 8'h00;
RAM[16'h6D19] = 8'h00;
RAM[16'h6D1A] = 8'h00;
RAM[16'h6D1B] = 8'h00;
RAM[16'h6D1C] = 8'h00;
RAM[16'h6D1D] = 8'h00;
RAM[16'h6D1E] = 8'h00;
RAM[16'h6D1F] = 8'h00;
RAM[16'h6D20] = 8'h00;
RAM[16'h6D21] = 8'h00;
RAM[16'h6D22] = 8'h00;
RAM[16'h6D23] = 8'h00;
RAM[16'h6D24] = 8'h00;
RAM[16'h6D25] = 8'h00;
RAM[16'h6D26] = 8'h00;
RAM[16'h6D27] = 8'h00;
RAM[16'h6D28] = 8'h00;
RAM[16'h6D29] = 8'h00;
RAM[16'h6D2A] = 8'h00;
RAM[16'h6D2B] = 8'h00;
RAM[16'h6D2C] = 8'h00;
RAM[16'h6D2D] = 8'h00;
RAM[16'h6D2E] = 8'h00;
RAM[16'h6D2F] = 8'h00;
RAM[16'h6D30] = 8'h00;
RAM[16'h6D31] = 8'h00;
RAM[16'h6D32] = 8'h00;
RAM[16'h6D33] = 8'h00;
RAM[16'h6D34] = 8'h00;
RAM[16'h6D35] = 8'h00;
RAM[16'h6D36] = 8'h00;
RAM[16'h6D37] = 8'h00;
RAM[16'h6D38] = 8'h00;
RAM[16'h6D39] = 8'h00;
RAM[16'h6D3A] = 8'h00;
RAM[16'h6D3B] = 8'h00;
RAM[16'h6D3C] = 8'h00;
RAM[16'h6D3D] = 8'h00;
RAM[16'h6D3E] = 8'h00;
RAM[16'h6D3F] = 8'h00;
RAM[16'h6D40] = 8'h00;
RAM[16'h6D41] = 8'h00;
RAM[16'h6D42] = 8'h00;
RAM[16'h6D43] = 8'h00;
RAM[16'h6D44] = 8'h00;
RAM[16'h6D45] = 8'h00;
RAM[16'h6D46] = 8'h00;
RAM[16'h6D47] = 8'h00;
RAM[16'h6D48] = 8'h00;
RAM[16'h6D49] = 8'h00;
RAM[16'h6D4A] = 8'h00;
RAM[16'h6D4B] = 8'h00;
RAM[16'h6D4C] = 8'h00;
RAM[16'h6D4D] = 8'h00;
RAM[16'h6D4E] = 8'h00;
RAM[16'h6D4F] = 8'h00;
RAM[16'h6D50] = 8'h00;
RAM[16'h6D51] = 8'h00;
RAM[16'h6D52] = 8'h00;
RAM[16'h6D53] = 8'h00;
RAM[16'h6D54] = 8'h00;
RAM[16'h6D55] = 8'h00;
RAM[16'h6D56] = 8'h00;
RAM[16'h6D57] = 8'h00;
RAM[16'h6D58] = 8'h00;
RAM[16'h6D59] = 8'h00;
RAM[16'h6D5A] = 8'h00;
RAM[16'h6D5B] = 8'h00;
RAM[16'h6D5C] = 8'h00;
RAM[16'h6D5D] = 8'h00;
RAM[16'h6D5E] = 8'h00;
RAM[16'h6D5F] = 8'h00;
RAM[16'h6D60] = 8'h00;
RAM[16'h6D61] = 8'h00;
RAM[16'h6D62] = 8'h00;
RAM[16'h6D63] = 8'h00;
RAM[16'h6D64] = 8'h00;
RAM[16'h6D65] = 8'h00;
RAM[16'h6D66] = 8'h00;
RAM[16'h6D67] = 8'h00;
RAM[16'h6D68] = 8'h00;
RAM[16'h6D69] = 8'h00;
RAM[16'h6D6A] = 8'h00;
RAM[16'h6D6B] = 8'h00;
RAM[16'h6D6C] = 8'h00;
RAM[16'h6D6D] = 8'h00;
RAM[16'h6D6E] = 8'h00;
RAM[16'h6D6F] = 8'h00;
RAM[16'h6D70] = 8'h00;
RAM[16'h6D71] = 8'h00;
RAM[16'h6D72] = 8'h00;
RAM[16'h6D73] = 8'h00;
RAM[16'h6D74] = 8'h00;
RAM[16'h6D75] = 8'h00;
RAM[16'h6D76] = 8'h00;
RAM[16'h6D77] = 8'h00;
RAM[16'h6D78] = 8'h00;
RAM[16'h6D79] = 8'h00;
RAM[16'h6D7A] = 8'h00;
RAM[16'h6D7B] = 8'h00;
RAM[16'h6D7C] = 8'h00;
RAM[16'h6D7D] = 8'h00;
RAM[16'h6D7E] = 8'h00;
RAM[16'h6D7F] = 8'h00;
RAM[16'h6D80] = 8'h00;
RAM[16'h6D81] = 8'h00;
RAM[16'h6D82] = 8'h00;
RAM[16'h6D83] = 8'h00;
RAM[16'h6D84] = 8'h00;
RAM[16'h6D85] = 8'h00;
RAM[16'h6D86] = 8'h00;
RAM[16'h6D87] = 8'h00;
RAM[16'h6D88] = 8'h00;
RAM[16'h6D89] = 8'h00;
RAM[16'h6D8A] = 8'h00;
RAM[16'h6D8B] = 8'h00;
RAM[16'h6D8C] = 8'h00;
RAM[16'h6D8D] = 8'h00;
RAM[16'h6D8E] = 8'h00;
RAM[16'h6D8F] = 8'h00;
RAM[16'h6D90] = 8'h00;
RAM[16'h6D91] = 8'h00;
RAM[16'h6D92] = 8'h00;
RAM[16'h6D93] = 8'h00;
RAM[16'h6D94] = 8'h00;
RAM[16'h6D95] = 8'h00;
RAM[16'h6D96] = 8'h00;
RAM[16'h6D97] = 8'h00;
RAM[16'h6D98] = 8'h00;
RAM[16'h6D99] = 8'h00;
RAM[16'h6D9A] = 8'h00;
RAM[16'h6D9B] = 8'h00;
RAM[16'h6D9C] = 8'h00;
RAM[16'h6D9D] = 8'h00;
RAM[16'h6D9E] = 8'h00;
RAM[16'h6D9F] = 8'h00;
RAM[16'h6DA0] = 8'h00;
RAM[16'h6DA1] = 8'h00;
RAM[16'h6DA2] = 8'h00;
RAM[16'h6DA3] = 8'h00;
RAM[16'h6DA4] = 8'h00;
RAM[16'h6DA5] = 8'h00;
RAM[16'h6DA6] = 8'h00;
RAM[16'h6DA7] = 8'h00;
RAM[16'h6DA8] = 8'h00;
RAM[16'h6DA9] = 8'h00;
RAM[16'h6DAA] = 8'h00;
RAM[16'h6DAB] = 8'h00;
RAM[16'h6DAC] = 8'h00;
RAM[16'h6DAD] = 8'h00;
RAM[16'h6DAE] = 8'h00;
RAM[16'h6DAF] = 8'h00;
RAM[16'h6DB0] = 8'h00;
RAM[16'h6DB1] = 8'h00;
RAM[16'h6DB2] = 8'h00;
RAM[16'h6DB3] = 8'h00;
RAM[16'h6DB4] = 8'h00;
RAM[16'h6DB5] = 8'h00;
RAM[16'h6DB6] = 8'h00;
RAM[16'h6DB7] = 8'h00;
RAM[16'h6DB8] = 8'h00;
RAM[16'h6DB9] = 8'h00;
RAM[16'h6DBA] = 8'h00;
RAM[16'h6DBB] = 8'h00;
RAM[16'h6DBC] = 8'h00;
RAM[16'h6DBD] = 8'h00;
RAM[16'h6DBE] = 8'h00;
RAM[16'h6DBF] = 8'h00;
RAM[16'h6DC0] = 8'h00;
RAM[16'h6DC1] = 8'h00;
RAM[16'h6DC2] = 8'h00;
RAM[16'h6DC3] = 8'h00;
RAM[16'h6DC4] = 8'h00;
RAM[16'h6DC5] = 8'h00;
RAM[16'h6DC6] = 8'h00;
RAM[16'h6DC7] = 8'h00;
RAM[16'h6DC8] = 8'h00;
RAM[16'h6DC9] = 8'h00;
RAM[16'h6DCA] = 8'h00;
RAM[16'h6DCB] = 8'h00;
RAM[16'h6DCC] = 8'h00;
RAM[16'h6DCD] = 8'h00;
RAM[16'h6DCE] = 8'h00;
RAM[16'h6DCF] = 8'h00;
RAM[16'h6DD0] = 8'h00;
RAM[16'h6DD1] = 8'h00;
RAM[16'h6DD2] = 8'h00;
RAM[16'h6DD3] = 8'h00;
RAM[16'h6DD4] = 8'h00;
RAM[16'h6DD5] = 8'h00;
RAM[16'h6DD6] = 8'h00;
RAM[16'h6DD7] = 8'h00;
RAM[16'h6DD8] = 8'h00;
RAM[16'h6DD9] = 8'h00;
RAM[16'h6DDA] = 8'h00;
RAM[16'h6DDB] = 8'h00;
RAM[16'h6DDC] = 8'h00;
RAM[16'h6DDD] = 8'h00;
RAM[16'h6DDE] = 8'h00;
RAM[16'h6DDF] = 8'h00;
RAM[16'h6DE0] = 8'h00;
RAM[16'h6DE1] = 8'h00;
RAM[16'h6DE2] = 8'h00;
RAM[16'h6DE3] = 8'h00;
RAM[16'h6DE4] = 8'h00;
RAM[16'h6DE5] = 8'h00;
RAM[16'h6DE6] = 8'h00;
RAM[16'h6DE7] = 8'h00;
RAM[16'h6DE8] = 8'h00;
RAM[16'h6DE9] = 8'h00;
RAM[16'h6DEA] = 8'h00;
RAM[16'h6DEB] = 8'h00;
RAM[16'h6DEC] = 8'h00;
RAM[16'h6DED] = 8'h00;
RAM[16'h6DEE] = 8'h00;
RAM[16'h6DEF] = 8'h00;
RAM[16'h6DF0] = 8'h00;
RAM[16'h6DF1] = 8'h00;
RAM[16'h6DF2] = 8'h00;
RAM[16'h6DF3] = 8'h00;
RAM[16'h6DF4] = 8'h00;
RAM[16'h6DF5] = 8'h00;
RAM[16'h6DF6] = 8'h00;
RAM[16'h6DF7] = 8'h00;
RAM[16'h6DF8] = 8'h00;
RAM[16'h6DF9] = 8'h00;
RAM[16'h6DFA] = 8'h00;
RAM[16'h6DFB] = 8'h00;
RAM[16'h6DFC] = 8'h00;
RAM[16'h6DFD] = 8'h00;
RAM[16'h6DFE] = 8'h00;
RAM[16'h6DFF] = 8'h00;
RAM[16'h6E00] = 8'h00;
RAM[16'h6E01] = 8'h00;
RAM[16'h6E02] = 8'h00;
RAM[16'h6E03] = 8'h00;
RAM[16'h6E04] = 8'h00;
RAM[16'h6E05] = 8'h00;
RAM[16'h6E06] = 8'h00;
RAM[16'h6E07] = 8'h00;
RAM[16'h6E08] = 8'h00;
RAM[16'h6E09] = 8'h00;
RAM[16'h6E0A] = 8'h00;
RAM[16'h6E0B] = 8'h00;
RAM[16'h6E0C] = 8'h00;
RAM[16'h6E0D] = 8'h00;
RAM[16'h6E0E] = 8'h00;
RAM[16'h6E0F] = 8'h00;
RAM[16'h6E10] = 8'h00;
RAM[16'h6E11] = 8'h00;
RAM[16'h6E12] = 8'h00;
RAM[16'h6E13] = 8'h00;
RAM[16'h6E14] = 8'h00;
RAM[16'h6E15] = 8'h00;
RAM[16'h6E16] = 8'h00;
RAM[16'h6E17] = 8'h00;
RAM[16'h6E18] = 8'h00;
RAM[16'h6E19] = 8'h00;
RAM[16'h6E1A] = 8'h00;
RAM[16'h6E1B] = 8'h00;
RAM[16'h6E1C] = 8'h00;
RAM[16'h6E1D] = 8'h00;
RAM[16'h6E1E] = 8'h00;
RAM[16'h6E1F] = 8'h00;
RAM[16'h6E20] = 8'h00;
RAM[16'h6E21] = 8'h00;
RAM[16'h6E22] = 8'h00;
RAM[16'h6E23] = 8'h00;
RAM[16'h6E24] = 8'h00;
RAM[16'h6E25] = 8'h00;
RAM[16'h6E26] = 8'h00;
RAM[16'h6E27] = 8'h00;
RAM[16'h6E28] = 8'h00;
RAM[16'h6E29] = 8'h00;
RAM[16'h6E2A] = 8'h00;
RAM[16'h6E2B] = 8'h00;
RAM[16'h6E2C] = 8'h00;
RAM[16'h6E2D] = 8'h00;
RAM[16'h6E2E] = 8'h00;
RAM[16'h6E2F] = 8'h00;
RAM[16'h6E30] = 8'h00;
RAM[16'h6E31] = 8'h00;
RAM[16'h6E32] = 8'h00;
RAM[16'h6E33] = 8'h00;
RAM[16'h6E34] = 8'h00;
RAM[16'h6E35] = 8'h00;
RAM[16'h6E36] = 8'h00;
RAM[16'h6E37] = 8'h00;
RAM[16'h6E38] = 8'h00;
RAM[16'h6E39] = 8'h00;
RAM[16'h6E3A] = 8'h00;
RAM[16'h6E3B] = 8'h00;
RAM[16'h6E3C] = 8'h00;
RAM[16'h6E3D] = 8'h00;
RAM[16'h6E3E] = 8'h00;
RAM[16'h6E3F] = 8'h00;
RAM[16'h6E40] = 8'h00;
RAM[16'h6E41] = 8'h00;
RAM[16'h6E42] = 8'h00;
RAM[16'h6E43] = 8'h00;
RAM[16'h6E44] = 8'h00;
RAM[16'h6E45] = 8'h00;
RAM[16'h6E46] = 8'h00;
RAM[16'h6E47] = 8'h00;
RAM[16'h6E48] = 8'h00;
RAM[16'h6E49] = 8'h00;
RAM[16'h6E4A] = 8'h00;
RAM[16'h6E4B] = 8'h00;
RAM[16'h6E4C] = 8'h00;
RAM[16'h6E4D] = 8'h00;
RAM[16'h6E4E] = 8'h00;
RAM[16'h6E4F] = 8'h00;
RAM[16'h6E50] = 8'h00;
RAM[16'h6E51] = 8'h00;
RAM[16'h6E52] = 8'h00;
RAM[16'h6E53] = 8'h00;
RAM[16'h6E54] = 8'h00;
RAM[16'h6E55] = 8'h00;
RAM[16'h6E56] = 8'h00;
RAM[16'h6E57] = 8'h00;
RAM[16'h6E58] = 8'h00;
RAM[16'h6E59] = 8'h00;
RAM[16'h6E5A] = 8'h00;
RAM[16'h6E5B] = 8'h00;
RAM[16'h6E5C] = 8'h00;
RAM[16'h6E5D] = 8'h00;
RAM[16'h6E5E] = 8'h00;
RAM[16'h6E5F] = 8'h00;
RAM[16'h6E60] = 8'h00;
RAM[16'h6E61] = 8'h00;
RAM[16'h6E62] = 8'h00;
RAM[16'h6E63] = 8'h00;
RAM[16'h6E64] = 8'h00;
RAM[16'h6E65] = 8'h00;
RAM[16'h6E66] = 8'h00;
RAM[16'h6E67] = 8'h00;
RAM[16'h6E68] = 8'h00;
RAM[16'h6E69] = 8'h00;
RAM[16'h6E6A] = 8'h00;
RAM[16'h6E6B] = 8'h00;
RAM[16'h6E6C] = 8'h00;
RAM[16'h6E6D] = 8'h00;
RAM[16'h6E6E] = 8'h00;
RAM[16'h6E6F] = 8'h00;
RAM[16'h6E70] = 8'h00;
RAM[16'h6E71] = 8'h00;
RAM[16'h6E72] = 8'h00;
RAM[16'h6E73] = 8'h00;
RAM[16'h6E74] = 8'h00;
RAM[16'h6E75] = 8'h00;
RAM[16'h6E76] = 8'h00;
RAM[16'h6E77] = 8'h00;
RAM[16'h6E78] = 8'h00;
RAM[16'h6E79] = 8'h00;
RAM[16'h6E7A] = 8'h00;
RAM[16'h6E7B] = 8'h00;
RAM[16'h6E7C] = 8'h00;
RAM[16'h6E7D] = 8'h00;
RAM[16'h6E7E] = 8'h00;
RAM[16'h6E7F] = 8'h00;
RAM[16'h6E80] = 8'h00;
RAM[16'h6E81] = 8'h00;
RAM[16'h6E82] = 8'h00;
RAM[16'h6E83] = 8'h00;
RAM[16'h6E84] = 8'h00;
RAM[16'h6E85] = 8'h00;
RAM[16'h6E86] = 8'h00;
RAM[16'h6E87] = 8'h00;
RAM[16'h6E88] = 8'h00;
RAM[16'h6E89] = 8'h00;
RAM[16'h6E8A] = 8'h00;
RAM[16'h6E8B] = 8'h00;
RAM[16'h6E8C] = 8'h00;
RAM[16'h6E8D] = 8'h00;
RAM[16'h6E8E] = 8'h00;
RAM[16'h6E8F] = 8'h00;
RAM[16'h6E90] = 8'h00;
RAM[16'h6E91] = 8'h00;
RAM[16'h6E92] = 8'h00;
RAM[16'h6E93] = 8'h00;
RAM[16'h6E94] = 8'h00;
RAM[16'h6E95] = 8'h00;
RAM[16'h6E96] = 8'h00;
RAM[16'h6E97] = 8'h00;
RAM[16'h6E98] = 8'h00;
RAM[16'h6E99] = 8'h00;
RAM[16'h6E9A] = 8'h00;
RAM[16'h6E9B] = 8'h00;
RAM[16'h6E9C] = 8'h00;
RAM[16'h6E9D] = 8'h00;
RAM[16'h6E9E] = 8'h00;
RAM[16'h6E9F] = 8'h00;
RAM[16'h6EA0] = 8'h00;
RAM[16'h6EA1] = 8'h00;
RAM[16'h6EA2] = 8'h00;
RAM[16'h6EA3] = 8'h00;
RAM[16'h6EA4] = 8'h00;
RAM[16'h6EA5] = 8'h00;
RAM[16'h6EA6] = 8'h00;
RAM[16'h6EA7] = 8'h00;
RAM[16'h6EA8] = 8'h00;
RAM[16'h6EA9] = 8'h00;
RAM[16'h6EAA] = 8'h00;
RAM[16'h6EAB] = 8'h00;
RAM[16'h6EAC] = 8'h00;
RAM[16'h6EAD] = 8'h00;
RAM[16'h6EAE] = 8'h00;
RAM[16'h6EAF] = 8'h00;
RAM[16'h6EB0] = 8'h00;
RAM[16'h6EB1] = 8'h00;
RAM[16'h6EB2] = 8'h00;
RAM[16'h6EB3] = 8'h00;
RAM[16'h6EB4] = 8'h00;
RAM[16'h6EB5] = 8'h00;
RAM[16'h6EB6] = 8'h00;
RAM[16'h6EB7] = 8'h00;
RAM[16'h6EB8] = 8'h00;
RAM[16'h6EB9] = 8'h00;
RAM[16'h6EBA] = 8'h00;
RAM[16'h6EBB] = 8'h00;
RAM[16'h6EBC] = 8'h00;
RAM[16'h6EBD] = 8'h00;
RAM[16'h6EBE] = 8'h00;
RAM[16'h6EBF] = 8'h00;
RAM[16'h6EC0] = 8'h00;
RAM[16'h6EC1] = 8'h00;
RAM[16'h6EC2] = 8'h00;
RAM[16'h6EC3] = 8'h00;
RAM[16'h6EC4] = 8'h00;
RAM[16'h6EC5] = 8'h00;
RAM[16'h6EC6] = 8'h00;
RAM[16'h6EC7] = 8'h00;
RAM[16'h6EC8] = 8'h00;
RAM[16'h6EC9] = 8'h00;
RAM[16'h6ECA] = 8'h00;
RAM[16'h6ECB] = 8'h00;
RAM[16'h6ECC] = 8'h00;
RAM[16'h6ECD] = 8'h00;
RAM[16'h6ECE] = 8'h00;
RAM[16'h6ECF] = 8'h00;
RAM[16'h6ED0] = 8'h00;
RAM[16'h6ED1] = 8'h00;
RAM[16'h6ED2] = 8'h00;
RAM[16'h6ED3] = 8'h00;
RAM[16'h6ED4] = 8'h00;
RAM[16'h6ED5] = 8'h00;
RAM[16'h6ED6] = 8'h00;
RAM[16'h6ED7] = 8'h00;
RAM[16'h6ED8] = 8'h00;
RAM[16'h6ED9] = 8'h00;
RAM[16'h6EDA] = 8'h00;
RAM[16'h6EDB] = 8'h00;
RAM[16'h6EDC] = 8'h00;
RAM[16'h6EDD] = 8'h00;
RAM[16'h6EDE] = 8'h00;
RAM[16'h6EDF] = 8'h00;
RAM[16'h6EE0] = 8'h00;
RAM[16'h6EE1] = 8'h00;
RAM[16'h6EE2] = 8'h00;
RAM[16'h6EE3] = 8'h00;
RAM[16'h6EE4] = 8'h00;
RAM[16'h6EE5] = 8'h00;
RAM[16'h6EE6] = 8'h00;
RAM[16'h6EE7] = 8'h00;
RAM[16'h6EE8] = 8'h00;
RAM[16'h6EE9] = 8'h00;
RAM[16'h6EEA] = 8'h00;
RAM[16'h6EEB] = 8'h00;
RAM[16'h6EEC] = 8'h00;
RAM[16'h6EED] = 8'h00;
RAM[16'h6EEE] = 8'h00;
RAM[16'h6EEF] = 8'h00;
RAM[16'h6EF0] = 8'h00;
RAM[16'h6EF1] = 8'h00;
RAM[16'h6EF2] = 8'h00;
RAM[16'h6EF3] = 8'h00;
RAM[16'h6EF4] = 8'h00;
RAM[16'h6EF5] = 8'h00;
RAM[16'h6EF6] = 8'h00;
RAM[16'h6EF7] = 8'h00;
RAM[16'h6EF8] = 8'h00;
RAM[16'h6EF9] = 8'h00;
RAM[16'h6EFA] = 8'h00;
RAM[16'h6EFB] = 8'h00;
RAM[16'h6EFC] = 8'h00;
RAM[16'h6EFD] = 8'h00;
RAM[16'h6EFE] = 8'h00;
RAM[16'h6EFF] = 8'h00;
RAM[16'h6F00] = 8'h00;
RAM[16'h6F01] = 8'h00;
RAM[16'h6F02] = 8'h00;
RAM[16'h6F03] = 8'h00;
RAM[16'h6F04] = 8'h00;
RAM[16'h6F05] = 8'h00;
RAM[16'h6F06] = 8'h00;
RAM[16'h6F07] = 8'h00;
RAM[16'h6F08] = 8'h00;
RAM[16'h6F09] = 8'h00;
RAM[16'h6F0A] = 8'h00;
RAM[16'h6F0B] = 8'h00;
RAM[16'h6F0C] = 8'h00;
RAM[16'h6F0D] = 8'h00;
RAM[16'h6F0E] = 8'h00;
RAM[16'h6F0F] = 8'h00;
RAM[16'h6F10] = 8'h00;
RAM[16'h6F11] = 8'h00;
RAM[16'h6F12] = 8'h00;
RAM[16'h6F13] = 8'h00;
RAM[16'h6F14] = 8'h00;
RAM[16'h6F15] = 8'h00;
RAM[16'h6F16] = 8'h00;
RAM[16'h6F17] = 8'h00;
RAM[16'h6F18] = 8'h00;
RAM[16'h6F19] = 8'h00;
RAM[16'h6F1A] = 8'h00;
RAM[16'h6F1B] = 8'h00;
RAM[16'h6F1C] = 8'h00;
RAM[16'h6F1D] = 8'h00;
RAM[16'h6F1E] = 8'h00;
RAM[16'h6F1F] = 8'h00;
RAM[16'h6F20] = 8'h00;
RAM[16'h6F21] = 8'h00;
RAM[16'h6F22] = 8'h00;
RAM[16'h6F23] = 8'h00;
RAM[16'h6F24] = 8'h00;
RAM[16'h6F25] = 8'h00;
RAM[16'h6F26] = 8'h00;
RAM[16'h6F27] = 8'h00;
RAM[16'h6F28] = 8'h00;
RAM[16'h6F29] = 8'h00;
RAM[16'h6F2A] = 8'h00;
RAM[16'h6F2B] = 8'h00;
RAM[16'h6F2C] = 8'h00;
RAM[16'h6F2D] = 8'h00;
RAM[16'h6F2E] = 8'h00;
RAM[16'h6F2F] = 8'h00;
RAM[16'h6F30] = 8'h00;
RAM[16'h6F31] = 8'h00;
RAM[16'h6F32] = 8'h00;
RAM[16'h6F33] = 8'h00;
RAM[16'h6F34] = 8'h00;
RAM[16'h6F35] = 8'h00;
RAM[16'h6F36] = 8'h00;
RAM[16'h6F37] = 8'h00;
RAM[16'h6F38] = 8'h00;
RAM[16'h6F39] = 8'h00;
RAM[16'h6F3A] = 8'h00;
RAM[16'h6F3B] = 8'h00;
RAM[16'h6F3C] = 8'h00;
RAM[16'h6F3D] = 8'h00;
RAM[16'h6F3E] = 8'h00;
RAM[16'h6F3F] = 8'h00;
RAM[16'h6F40] = 8'h00;
RAM[16'h6F41] = 8'h00;
RAM[16'h6F42] = 8'h00;
RAM[16'h6F43] = 8'h00;
RAM[16'h6F44] = 8'h00;
RAM[16'h6F45] = 8'h00;
RAM[16'h6F46] = 8'h00;
RAM[16'h6F47] = 8'h00;
RAM[16'h6F48] = 8'h00;
RAM[16'h6F49] = 8'h00;
RAM[16'h6F4A] = 8'h00;
RAM[16'h6F4B] = 8'h00;
RAM[16'h6F4C] = 8'h00;
RAM[16'h6F4D] = 8'h00;
RAM[16'h6F4E] = 8'h00;
RAM[16'h6F4F] = 8'h00;
RAM[16'h6F50] = 8'h00;
RAM[16'h6F51] = 8'h00;
RAM[16'h6F52] = 8'h00;
RAM[16'h6F53] = 8'h00;
RAM[16'h6F54] = 8'h00;
RAM[16'h6F55] = 8'h00;
RAM[16'h6F56] = 8'h00;
RAM[16'h6F57] = 8'h00;
RAM[16'h6F58] = 8'h00;
RAM[16'h6F59] = 8'h00;
RAM[16'h6F5A] = 8'h00;
RAM[16'h6F5B] = 8'h00;
RAM[16'h6F5C] = 8'h00;
RAM[16'h6F5D] = 8'h00;
RAM[16'h6F5E] = 8'h00;
RAM[16'h6F5F] = 8'h00;
RAM[16'h6F60] = 8'h00;
RAM[16'h6F61] = 8'h00;
RAM[16'h6F62] = 8'h00;
RAM[16'h6F63] = 8'h00;
RAM[16'h6F64] = 8'h00;
RAM[16'h6F65] = 8'h00;
RAM[16'h6F66] = 8'h00;
RAM[16'h6F67] = 8'h00;
RAM[16'h6F68] = 8'h00;
RAM[16'h6F69] = 8'h00;
RAM[16'h6F6A] = 8'h00;
RAM[16'h6F6B] = 8'h00;
RAM[16'h6F6C] = 8'h00;
RAM[16'h6F6D] = 8'h00;
RAM[16'h6F6E] = 8'h00;
RAM[16'h6F6F] = 8'h00;
RAM[16'h6F70] = 8'h00;
RAM[16'h6F71] = 8'h00;
RAM[16'h6F72] = 8'h00;
RAM[16'h6F73] = 8'h00;
RAM[16'h6F74] = 8'h00;
RAM[16'h6F75] = 8'h00;
RAM[16'h6F76] = 8'h00;
RAM[16'h6F77] = 8'h00;
RAM[16'h6F78] = 8'h00;
RAM[16'h6F79] = 8'h00;
RAM[16'h6F7A] = 8'h00;
RAM[16'h6F7B] = 8'h00;
RAM[16'h6F7C] = 8'h00;
RAM[16'h6F7D] = 8'h00;
RAM[16'h6F7E] = 8'h00;
RAM[16'h6F7F] = 8'h00;
RAM[16'h6F80] = 8'h00;
RAM[16'h6F81] = 8'h00;
RAM[16'h6F82] = 8'h00;
RAM[16'h6F83] = 8'h00;
RAM[16'h6F84] = 8'h00;
RAM[16'h6F85] = 8'h00;
RAM[16'h6F86] = 8'h00;
RAM[16'h6F87] = 8'h00;
RAM[16'h6F88] = 8'h00;
RAM[16'h6F89] = 8'h00;
RAM[16'h6F8A] = 8'h00;
RAM[16'h6F8B] = 8'h00;
RAM[16'h6F8C] = 8'h00;
RAM[16'h6F8D] = 8'h00;
RAM[16'h6F8E] = 8'h00;
RAM[16'h6F8F] = 8'h00;
RAM[16'h6F90] = 8'h00;
RAM[16'h6F91] = 8'h00;
RAM[16'h6F92] = 8'h00;
RAM[16'h6F93] = 8'h00;
RAM[16'h6F94] = 8'h00;
RAM[16'h6F95] = 8'h00;
RAM[16'h6F96] = 8'h00;
RAM[16'h6F97] = 8'h00;
RAM[16'h6F98] = 8'h00;
RAM[16'h6F99] = 8'h00;
RAM[16'h6F9A] = 8'h00;
RAM[16'h6F9B] = 8'h00;
RAM[16'h6F9C] = 8'h00;
RAM[16'h6F9D] = 8'h00;
RAM[16'h6F9E] = 8'h00;
RAM[16'h6F9F] = 8'h00;
RAM[16'h6FA0] = 8'h00;
RAM[16'h6FA1] = 8'h00;
RAM[16'h6FA2] = 8'h00;
RAM[16'h6FA3] = 8'h00;
RAM[16'h6FA4] = 8'h00;
RAM[16'h6FA5] = 8'h00;
RAM[16'h6FA6] = 8'h00;
RAM[16'h6FA7] = 8'h00;
RAM[16'h6FA8] = 8'h00;
RAM[16'h6FA9] = 8'h00;
RAM[16'h6FAA] = 8'h00;
RAM[16'h6FAB] = 8'h00;
RAM[16'h6FAC] = 8'h00;
RAM[16'h6FAD] = 8'h00;
RAM[16'h6FAE] = 8'h00;
RAM[16'h6FAF] = 8'h00;
RAM[16'h6FB0] = 8'h00;
RAM[16'h6FB1] = 8'h00;
RAM[16'h6FB2] = 8'h00;
RAM[16'h6FB3] = 8'h00;
RAM[16'h6FB4] = 8'h00;
RAM[16'h6FB5] = 8'h00;
RAM[16'h6FB6] = 8'h00;
RAM[16'h6FB7] = 8'h00;
RAM[16'h6FB8] = 8'h00;
RAM[16'h6FB9] = 8'h00;
RAM[16'h6FBA] = 8'h00;
RAM[16'h6FBB] = 8'h00;
RAM[16'h6FBC] = 8'h00;
RAM[16'h6FBD] = 8'h00;
RAM[16'h6FBE] = 8'h00;
RAM[16'h6FBF] = 8'h00;
RAM[16'h6FC0] = 8'h00;
RAM[16'h6FC1] = 8'h00;
RAM[16'h6FC2] = 8'h00;
RAM[16'h6FC3] = 8'h00;
RAM[16'h6FC4] = 8'h00;
RAM[16'h6FC5] = 8'h00;
RAM[16'h6FC6] = 8'h00;
RAM[16'h6FC7] = 8'h00;
RAM[16'h6FC8] = 8'h00;
RAM[16'h6FC9] = 8'h00;
RAM[16'h6FCA] = 8'h00;
RAM[16'h6FCB] = 8'h00;
RAM[16'h6FCC] = 8'h00;
RAM[16'h6FCD] = 8'h00;
RAM[16'h6FCE] = 8'h00;
RAM[16'h6FCF] = 8'h00;
RAM[16'h6FD0] = 8'h00;
RAM[16'h6FD1] = 8'h00;
RAM[16'h6FD2] = 8'h00;
RAM[16'h6FD3] = 8'h00;
RAM[16'h6FD4] = 8'h00;
RAM[16'h6FD5] = 8'h00;
RAM[16'h6FD6] = 8'h00;
RAM[16'h6FD7] = 8'h00;
RAM[16'h6FD8] = 8'h00;
RAM[16'h6FD9] = 8'h00;
RAM[16'h6FDA] = 8'h00;
RAM[16'h6FDB] = 8'h00;
RAM[16'h6FDC] = 8'h00;
RAM[16'h6FDD] = 8'h00;
RAM[16'h6FDE] = 8'h00;
RAM[16'h6FDF] = 8'h00;
RAM[16'h6FE0] = 8'h00;
RAM[16'h6FE1] = 8'h00;
RAM[16'h6FE2] = 8'h00;
RAM[16'h6FE3] = 8'h00;
RAM[16'h6FE4] = 8'h00;
RAM[16'h6FE5] = 8'h00;
RAM[16'h6FE6] = 8'h00;
RAM[16'h6FE7] = 8'h00;
RAM[16'h6FE8] = 8'h00;
RAM[16'h6FE9] = 8'h00;
RAM[16'h6FEA] = 8'h00;
RAM[16'h6FEB] = 8'h00;
RAM[16'h6FEC] = 8'h00;
RAM[16'h6FED] = 8'h00;
RAM[16'h6FEE] = 8'h00;
RAM[16'h6FEF] = 8'h00;
RAM[16'h6FF0] = 8'h00;
RAM[16'h6FF1] = 8'h00;
RAM[16'h6FF2] = 8'h00;
RAM[16'h6FF3] = 8'h00;
RAM[16'h6FF4] = 8'h00;
RAM[16'h6FF5] = 8'h00;
RAM[16'h6FF6] = 8'h00;
RAM[16'h6FF7] = 8'h00;
RAM[16'h6FF8] = 8'h00;
RAM[16'h6FF9] = 8'h00;
RAM[16'h6FFA] = 8'h00;
RAM[16'h6FFB] = 8'h00;
RAM[16'h6FFC] = 8'h00;
RAM[16'h6FFD] = 8'h00;
RAM[16'h6FFE] = 8'h00;
RAM[16'h6FFF] = 8'h00;
RAM[16'h7000] = 8'h00;
RAM[16'h7001] = 8'h00;
RAM[16'h7002] = 8'h00;
RAM[16'h7003] = 8'h00;
RAM[16'h7004] = 8'h00;
RAM[16'h7005] = 8'h00;
RAM[16'h7006] = 8'h00;
RAM[16'h7007] = 8'h00;
RAM[16'h7008] = 8'h00;
RAM[16'h7009] = 8'h00;
RAM[16'h700A] = 8'h00;
RAM[16'h700B] = 8'h00;
RAM[16'h700C] = 8'h00;
RAM[16'h700D] = 8'h00;
RAM[16'h700E] = 8'h00;
RAM[16'h700F] = 8'h00;
RAM[16'h7010] = 8'h00;
RAM[16'h7011] = 8'h00;
RAM[16'h7012] = 8'h00;
RAM[16'h7013] = 8'h00;
RAM[16'h7014] = 8'h00;
RAM[16'h7015] = 8'h00;
RAM[16'h7016] = 8'h00;
RAM[16'h7017] = 8'h00;
RAM[16'h7018] = 8'h00;
RAM[16'h7019] = 8'h00;
RAM[16'h701A] = 8'h00;
RAM[16'h701B] = 8'h00;
RAM[16'h701C] = 8'h00;
RAM[16'h701D] = 8'h00;
RAM[16'h701E] = 8'h00;
RAM[16'h701F] = 8'h00;
RAM[16'h7020] = 8'h00;
RAM[16'h7021] = 8'h00;
RAM[16'h7022] = 8'h00;
RAM[16'h7023] = 8'h00;
RAM[16'h7024] = 8'h00;
RAM[16'h7025] = 8'h00;
RAM[16'h7026] = 8'h00;
RAM[16'h7027] = 8'h00;
RAM[16'h7028] = 8'h00;
RAM[16'h7029] = 8'h00;
RAM[16'h702A] = 8'h00;
RAM[16'h702B] = 8'h00;
RAM[16'h702C] = 8'h00;
RAM[16'h702D] = 8'h00;
RAM[16'h702E] = 8'h00;
RAM[16'h702F] = 8'h00;
RAM[16'h7030] = 8'h00;
RAM[16'h7031] = 8'h00;
RAM[16'h7032] = 8'h00;
RAM[16'h7033] = 8'h00;
RAM[16'h7034] = 8'h00;
RAM[16'h7035] = 8'h00;
RAM[16'h7036] = 8'h00;
RAM[16'h7037] = 8'h00;
RAM[16'h7038] = 8'h00;
RAM[16'h7039] = 8'h00;
RAM[16'h703A] = 8'h00;
RAM[16'h703B] = 8'h00;
RAM[16'h703C] = 8'h00;
RAM[16'h703D] = 8'h00;
RAM[16'h703E] = 8'h00;
RAM[16'h703F] = 8'h00;
RAM[16'h7040] = 8'h00;
RAM[16'h7041] = 8'h00;
RAM[16'h7042] = 8'h00;
RAM[16'h7043] = 8'h00;
RAM[16'h7044] = 8'h00;
RAM[16'h7045] = 8'h00;
RAM[16'h7046] = 8'h00;
RAM[16'h7047] = 8'h00;
RAM[16'h7048] = 8'h00;
RAM[16'h7049] = 8'h00;
RAM[16'h704A] = 8'h00;
RAM[16'h704B] = 8'h00;
RAM[16'h704C] = 8'h00;
RAM[16'h704D] = 8'h00;
RAM[16'h704E] = 8'h00;
RAM[16'h704F] = 8'h00;
RAM[16'h7050] = 8'h00;
RAM[16'h7051] = 8'h00;
RAM[16'h7052] = 8'h00;
RAM[16'h7053] = 8'h00;
RAM[16'h7054] = 8'h00;
RAM[16'h7055] = 8'h00;
RAM[16'h7056] = 8'h00;
RAM[16'h7057] = 8'h00;
RAM[16'h7058] = 8'h00;
RAM[16'h7059] = 8'h00;
RAM[16'h705A] = 8'h00;
RAM[16'h705B] = 8'h00;
RAM[16'h705C] = 8'h00;
RAM[16'h705D] = 8'h00;
RAM[16'h705E] = 8'h00;
RAM[16'h705F] = 8'h00;
RAM[16'h7060] = 8'h00;
RAM[16'h7061] = 8'h00;
RAM[16'h7062] = 8'h00;
RAM[16'h7063] = 8'h00;
RAM[16'h7064] = 8'h00;
RAM[16'h7065] = 8'h00;
RAM[16'h7066] = 8'h00;
RAM[16'h7067] = 8'h00;
RAM[16'h7068] = 8'h00;
RAM[16'h7069] = 8'h00;
RAM[16'h706A] = 8'h00;
RAM[16'h706B] = 8'h00;
RAM[16'h706C] = 8'h00;
RAM[16'h706D] = 8'h00;
RAM[16'h706E] = 8'h00;
RAM[16'h706F] = 8'h00;
RAM[16'h7070] = 8'h00;
RAM[16'h7071] = 8'h00;
RAM[16'h7072] = 8'h00;
RAM[16'h7073] = 8'h00;
RAM[16'h7074] = 8'h00;
RAM[16'h7075] = 8'h00;
RAM[16'h7076] = 8'h00;
RAM[16'h7077] = 8'h00;
RAM[16'h7078] = 8'h00;
RAM[16'h7079] = 8'h00;
RAM[16'h707A] = 8'h00;
RAM[16'h707B] = 8'h00;
RAM[16'h707C] = 8'h00;
RAM[16'h707D] = 8'h00;
RAM[16'h707E] = 8'h00;
RAM[16'h707F] = 8'h00;
RAM[16'h7080] = 8'h00;
RAM[16'h7081] = 8'h00;
RAM[16'h7082] = 8'h00;
RAM[16'h7083] = 8'h00;
RAM[16'h7084] = 8'h00;
RAM[16'h7085] = 8'h00;
RAM[16'h7086] = 8'h00;
RAM[16'h7087] = 8'h00;
RAM[16'h7088] = 8'h00;
RAM[16'h7089] = 8'h00;
RAM[16'h708A] = 8'h00;
RAM[16'h708B] = 8'h00;
RAM[16'h708C] = 8'h00;
RAM[16'h708D] = 8'h00;
RAM[16'h708E] = 8'h00;
RAM[16'h708F] = 8'h00;
RAM[16'h7090] = 8'h00;
RAM[16'h7091] = 8'h00;
RAM[16'h7092] = 8'h00;
RAM[16'h7093] = 8'h00;
RAM[16'h7094] = 8'h00;
RAM[16'h7095] = 8'h00;
RAM[16'h7096] = 8'h00;
RAM[16'h7097] = 8'h00;
RAM[16'h7098] = 8'h00;
RAM[16'h7099] = 8'h00;
RAM[16'h709A] = 8'h00;
RAM[16'h709B] = 8'h00;
RAM[16'h709C] = 8'h00;
RAM[16'h709D] = 8'h00;
RAM[16'h709E] = 8'h00;
RAM[16'h709F] = 8'h00;
RAM[16'h70A0] = 8'h00;
RAM[16'h70A1] = 8'h00;
RAM[16'h70A2] = 8'h00;
RAM[16'h70A3] = 8'h00;
RAM[16'h70A4] = 8'h00;
RAM[16'h70A5] = 8'h00;
RAM[16'h70A6] = 8'h00;
RAM[16'h70A7] = 8'h00;
RAM[16'h70A8] = 8'h00;
RAM[16'h70A9] = 8'h00;
RAM[16'h70AA] = 8'h00;
RAM[16'h70AB] = 8'h00;
RAM[16'h70AC] = 8'h00;
RAM[16'h70AD] = 8'h00;
RAM[16'h70AE] = 8'h00;
RAM[16'h70AF] = 8'h00;
RAM[16'h70B0] = 8'h00;
RAM[16'h70B1] = 8'h00;
RAM[16'h70B2] = 8'h00;
RAM[16'h70B3] = 8'h00;
RAM[16'h70B4] = 8'h00;
RAM[16'h70B5] = 8'h00;
RAM[16'h70B6] = 8'h00;
RAM[16'h70B7] = 8'h00;
RAM[16'h70B8] = 8'h00;
RAM[16'h70B9] = 8'h00;
RAM[16'h70BA] = 8'h00;
RAM[16'h70BB] = 8'h00;
RAM[16'h70BC] = 8'h00;
RAM[16'h70BD] = 8'h00;
RAM[16'h70BE] = 8'h00;
RAM[16'h70BF] = 8'h00;
RAM[16'h70C0] = 8'h00;
RAM[16'h70C1] = 8'h00;
RAM[16'h70C2] = 8'h00;
RAM[16'h70C3] = 8'h00;
RAM[16'h70C4] = 8'h00;
RAM[16'h70C5] = 8'h00;
RAM[16'h70C6] = 8'h00;
RAM[16'h70C7] = 8'h00;
RAM[16'h70C8] = 8'h00;
RAM[16'h70C9] = 8'h00;
RAM[16'h70CA] = 8'h00;
RAM[16'h70CB] = 8'h00;
RAM[16'h70CC] = 8'h00;
RAM[16'h70CD] = 8'h00;
RAM[16'h70CE] = 8'h00;
RAM[16'h70CF] = 8'h00;
RAM[16'h70D0] = 8'h00;
RAM[16'h70D1] = 8'h00;
RAM[16'h70D2] = 8'h00;
RAM[16'h70D3] = 8'h00;
RAM[16'h70D4] = 8'h00;
RAM[16'h70D5] = 8'h00;
RAM[16'h70D6] = 8'h00;
RAM[16'h70D7] = 8'h00;
RAM[16'h70D8] = 8'h00;
RAM[16'h70D9] = 8'h00;
RAM[16'h70DA] = 8'h00;
RAM[16'h70DB] = 8'h00;
RAM[16'h70DC] = 8'h00;
RAM[16'h70DD] = 8'h00;
RAM[16'h70DE] = 8'h00;
RAM[16'h70DF] = 8'h00;
RAM[16'h70E0] = 8'h00;
RAM[16'h70E1] = 8'h00;
RAM[16'h70E2] = 8'h00;
RAM[16'h70E3] = 8'h00;
RAM[16'h70E4] = 8'h00;
RAM[16'h70E5] = 8'h00;
RAM[16'h70E6] = 8'h00;
RAM[16'h70E7] = 8'h00;
RAM[16'h70E8] = 8'h00;
RAM[16'h70E9] = 8'h00;
RAM[16'h70EA] = 8'h00;
RAM[16'h70EB] = 8'h00;
RAM[16'h70EC] = 8'h00;
RAM[16'h70ED] = 8'h00;
RAM[16'h70EE] = 8'h00;
RAM[16'h70EF] = 8'h00;
RAM[16'h70F0] = 8'h00;
RAM[16'h70F1] = 8'h00;
RAM[16'h70F2] = 8'h00;
RAM[16'h70F3] = 8'h00;
RAM[16'h70F4] = 8'h00;
RAM[16'h70F5] = 8'h00;
RAM[16'h70F6] = 8'h00;
RAM[16'h70F7] = 8'h00;
RAM[16'h70F8] = 8'h00;
RAM[16'h70F9] = 8'h00;
RAM[16'h70FA] = 8'h00;
RAM[16'h70FB] = 8'h00;
RAM[16'h70FC] = 8'h00;
RAM[16'h70FD] = 8'h00;
RAM[16'h70FE] = 8'h00;
RAM[16'h70FF] = 8'h00;
RAM[16'h7100] = 8'h00;
RAM[16'h7101] = 8'h00;
RAM[16'h7102] = 8'h00;
RAM[16'h7103] = 8'h00;
RAM[16'h7104] = 8'h00;
RAM[16'h7105] = 8'h00;
RAM[16'h7106] = 8'h00;
RAM[16'h7107] = 8'h00;
RAM[16'h7108] = 8'h00;
RAM[16'h7109] = 8'h00;
RAM[16'h710A] = 8'h00;
RAM[16'h710B] = 8'h00;
RAM[16'h710C] = 8'h00;
RAM[16'h710D] = 8'h00;
RAM[16'h710E] = 8'h00;
RAM[16'h710F] = 8'h00;
RAM[16'h7110] = 8'h00;
RAM[16'h7111] = 8'h00;
RAM[16'h7112] = 8'h00;
RAM[16'h7113] = 8'h00;
RAM[16'h7114] = 8'h00;
RAM[16'h7115] = 8'h00;
RAM[16'h7116] = 8'h00;
RAM[16'h7117] = 8'h00;
RAM[16'h7118] = 8'h00;
RAM[16'h7119] = 8'h00;
RAM[16'h711A] = 8'h00;
RAM[16'h711B] = 8'h00;
RAM[16'h711C] = 8'h00;
RAM[16'h711D] = 8'h00;
RAM[16'h711E] = 8'h00;
RAM[16'h711F] = 8'h00;
RAM[16'h7120] = 8'h00;
RAM[16'h7121] = 8'h00;
RAM[16'h7122] = 8'h00;
RAM[16'h7123] = 8'h00;
RAM[16'h7124] = 8'h00;
RAM[16'h7125] = 8'h00;
RAM[16'h7126] = 8'h00;
RAM[16'h7127] = 8'h00;
RAM[16'h7128] = 8'h00;
RAM[16'h7129] = 8'h00;
RAM[16'h712A] = 8'h00;
RAM[16'h712B] = 8'h00;
RAM[16'h712C] = 8'h00;
RAM[16'h712D] = 8'h00;
RAM[16'h712E] = 8'h00;
RAM[16'h712F] = 8'h00;
RAM[16'h7130] = 8'h00;
RAM[16'h7131] = 8'h00;
RAM[16'h7132] = 8'h00;
RAM[16'h7133] = 8'h00;
RAM[16'h7134] = 8'h00;
RAM[16'h7135] = 8'h00;
RAM[16'h7136] = 8'h00;
RAM[16'h7137] = 8'h00;
RAM[16'h7138] = 8'h00;
RAM[16'h7139] = 8'h00;
RAM[16'h713A] = 8'h00;
RAM[16'h713B] = 8'h00;
RAM[16'h713C] = 8'h00;
RAM[16'h713D] = 8'h00;
RAM[16'h713E] = 8'h00;
RAM[16'h713F] = 8'h00;
RAM[16'h7140] = 8'h00;
RAM[16'h7141] = 8'h00;
RAM[16'h7142] = 8'h00;
RAM[16'h7143] = 8'h00;
RAM[16'h7144] = 8'h00;
RAM[16'h7145] = 8'h00;
RAM[16'h7146] = 8'h00;
RAM[16'h7147] = 8'h00;
RAM[16'h7148] = 8'h00;
RAM[16'h7149] = 8'h00;
RAM[16'h714A] = 8'h00;
RAM[16'h714B] = 8'h00;
RAM[16'h714C] = 8'h00;
RAM[16'h714D] = 8'h00;
RAM[16'h714E] = 8'h00;
RAM[16'h714F] = 8'h00;
RAM[16'h7150] = 8'h00;
RAM[16'h7151] = 8'h00;
RAM[16'h7152] = 8'h00;
RAM[16'h7153] = 8'h00;
RAM[16'h7154] = 8'h00;
RAM[16'h7155] = 8'h00;
RAM[16'h7156] = 8'h00;
RAM[16'h7157] = 8'h00;
RAM[16'h7158] = 8'h00;
RAM[16'h7159] = 8'h00;
RAM[16'h715A] = 8'h00;
RAM[16'h715B] = 8'h00;
RAM[16'h715C] = 8'h00;
RAM[16'h715D] = 8'h00;
RAM[16'h715E] = 8'h00;
RAM[16'h715F] = 8'h00;
RAM[16'h7160] = 8'h00;
RAM[16'h7161] = 8'h00;
RAM[16'h7162] = 8'h00;
RAM[16'h7163] = 8'h00;
RAM[16'h7164] = 8'h00;
RAM[16'h7165] = 8'h00;
RAM[16'h7166] = 8'h00;
RAM[16'h7167] = 8'h00;
RAM[16'h7168] = 8'h00;
RAM[16'h7169] = 8'h00;
RAM[16'h716A] = 8'h00;
RAM[16'h716B] = 8'h00;
RAM[16'h716C] = 8'h00;
RAM[16'h716D] = 8'h00;
RAM[16'h716E] = 8'h00;
RAM[16'h716F] = 8'h00;
RAM[16'h7170] = 8'h00;
RAM[16'h7171] = 8'h00;
RAM[16'h7172] = 8'h00;
RAM[16'h7173] = 8'h00;
RAM[16'h7174] = 8'h00;
RAM[16'h7175] = 8'h00;
RAM[16'h7176] = 8'h00;
RAM[16'h7177] = 8'h00;
RAM[16'h7178] = 8'h00;
RAM[16'h7179] = 8'h00;
RAM[16'h717A] = 8'h00;
RAM[16'h717B] = 8'h00;
RAM[16'h717C] = 8'h00;
RAM[16'h717D] = 8'h00;
RAM[16'h717E] = 8'h00;
RAM[16'h717F] = 8'h00;
RAM[16'h7180] = 8'h00;
RAM[16'h7181] = 8'h00;
RAM[16'h7182] = 8'h00;
RAM[16'h7183] = 8'h00;
RAM[16'h7184] = 8'h00;
RAM[16'h7185] = 8'h00;
RAM[16'h7186] = 8'h00;
RAM[16'h7187] = 8'h00;
RAM[16'h7188] = 8'h00;
RAM[16'h7189] = 8'h00;
RAM[16'h718A] = 8'h00;
RAM[16'h718B] = 8'h00;
RAM[16'h718C] = 8'h00;
RAM[16'h718D] = 8'h00;
RAM[16'h718E] = 8'h00;
RAM[16'h718F] = 8'h00;
RAM[16'h7190] = 8'h00;
RAM[16'h7191] = 8'h00;
RAM[16'h7192] = 8'h00;
RAM[16'h7193] = 8'h00;
RAM[16'h7194] = 8'h00;
RAM[16'h7195] = 8'h00;
RAM[16'h7196] = 8'h00;
RAM[16'h7197] = 8'h00;
RAM[16'h7198] = 8'h00;
RAM[16'h7199] = 8'h00;
RAM[16'h719A] = 8'h00;
RAM[16'h719B] = 8'h00;
RAM[16'h719C] = 8'h00;
RAM[16'h719D] = 8'h00;
RAM[16'h719E] = 8'h00;
RAM[16'h719F] = 8'h00;
RAM[16'h71A0] = 8'h00;
RAM[16'h71A1] = 8'h00;
RAM[16'h71A2] = 8'h00;
RAM[16'h71A3] = 8'h00;
RAM[16'h71A4] = 8'h00;
RAM[16'h71A5] = 8'h00;
RAM[16'h71A6] = 8'h00;
RAM[16'h71A7] = 8'h00;
RAM[16'h71A8] = 8'h00;
RAM[16'h71A9] = 8'h00;
RAM[16'h71AA] = 8'h00;
RAM[16'h71AB] = 8'h00;
RAM[16'h71AC] = 8'h00;
RAM[16'h71AD] = 8'h00;
RAM[16'h71AE] = 8'h00;
RAM[16'h71AF] = 8'h00;
RAM[16'h71B0] = 8'h00;
RAM[16'h71B1] = 8'h00;
RAM[16'h71B2] = 8'h00;
RAM[16'h71B3] = 8'h00;
RAM[16'h71B4] = 8'h00;
RAM[16'h71B5] = 8'h00;
RAM[16'h71B6] = 8'h00;
RAM[16'h71B7] = 8'h00;
RAM[16'h71B8] = 8'h00;
RAM[16'h71B9] = 8'h00;
RAM[16'h71BA] = 8'h00;
RAM[16'h71BB] = 8'h00;
RAM[16'h71BC] = 8'h00;
RAM[16'h71BD] = 8'h00;
RAM[16'h71BE] = 8'h00;
RAM[16'h71BF] = 8'h00;
RAM[16'h71C0] = 8'h00;
RAM[16'h71C1] = 8'h00;
RAM[16'h71C2] = 8'h00;
RAM[16'h71C3] = 8'h00;
RAM[16'h71C4] = 8'h00;
RAM[16'h71C5] = 8'h00;
RAM[16'h71C6] = 8'h00;
RAM[16'h71C7] = 8'h00;
RAM[16'h71C8] = 8'h00;
RAM[16'h71C9] = 8'h00;
RAM[16'h71CA] = 8'h00;
RAM[16'h71CB] = 8'h00;
RAM[16'h71CC] = 8'h00;
RAM[16'h71CD] = 8'h00;
RAM[16'h71CE] = 8'h00;
RAM[16'h71CF] = 8'h00;
RAM[16'h71D0] = 8'h00;
RAM[16'h71D1] = 8'h00;
RAM[16'h71D2] = 8'h00;
RAM[16'h71D3] = 8'h00;
RAM[16'h71D4] = 8'h00;
RAM[16'h71D5] = 8'h00;
RAM[16'h71D6] = 8'h00;
RAM[16'h71D7] = 8'h00;
RAM[16'h71D8] = 8'h00;
RAM[16'h71D9] = 8'h00;
RAM[16'h71DA] = 8'h00;
RAM[16'h71DB] = 8'h00;
RAM[16'h71DC] = 8'h00;
RAM[16'h71DD] = 8'h00;
RAM[16'h71DE] = 8'h00;
RAM[16'h71DF] = 8'h00;
RAM[16'h71E0] = 8'h00;
RAM[16'h71E1] = 8'h00;
RAM[16'h71E2] = 8'h00;
RAM[16'h71E3] = 8'h00;
RAM[16'h71E4] = 8'h00;
RAM[16'h71E5] = 8'h00;
RAM[16'h71E6] = 8'h00;
RAM[16'h71E7] = 8'h00;
RAM[16'h71E8] = 8'h00;
RAM[16'h71E9] = 8'h00;
RAM[16'h71EA] = 8'h00;
RAM[16'h71EB] = 8'h00;
RAM[16'h71EC] = 8'h00;
RAM[16'h71ED] = 8'h00;
RAM[16'h71EE] = 8'h00;
RAM[16'h71EF] = 8'h00;
RAM[16'h71F0] = 8'h00;
RAM[16'h71F1] = 8'h00;
RAM[16'h71F2] = 8'h00;
RAM[16'h71F3] = 8'h00;
RAM[16'h71F4] = 8'h00;
RAM[16'h71F5] = 8'h00;
RAM[16'h71F6] = 8'h00;
RAM[16'h71F7] = 8'h00;
RAM[16'h71F8] = 8'h00;
RAM[16'h71F9] = 8'h00;
RAM[16'h71FA] = 8'h00;
RAM[16'h71FB] = 8'h00;
RAM[16'h71FC] = 8'h00;
RAM[16'h71FD] = 8'h00;
RAM[16'h71FE] = 8'h00;
RAM[16'h71FF] = 8'h00;
RAM[16'h7200] = 8'h00;
RAM[16'h7201] = 8'h00;
RAM[16'h7202] = 8'h00;
RAM[16'h7203] = 8'h00;
RAM[16'h7204] = 8'h00;
RAM[16'h7205] = 8'h00;
RAM[16'h7206] = 8'h00;
RAM[16'h7207] = 8'h00;
RAM[16'h7208] = 8'h00;
RAM[16'h7209] = 8'h00;
RAM[16'h720A] = 8'h00;
RAM[16'h720B] = 8'h00;
RAM[16'h720C] = 8'h00;
RAM[16'h720D] = 8'h00;
RAM[16'h720E] = 8'h00;
RAM[16'h720F] = 8'h00;
RAM[16'h7210] = 8'h00;
RAM[16'h7211] = 8'h00;
RAM[16'h7212] = 8'h00;
RAM[16'h7213] = 8'h00;
RAM[16'h7214] = 8'h00;
RAM[16'h7215] = 8'h00;
RAM[16'h7216] = 8'h00;
RAM[16'h7217] = 8'h00;
RAM[16'h7218] = 8'h00;
RAM[16'h7219] = 8'h00;
RAM[16'h721A] = 8'h00;
RAM[16'h721B] = 8'h00;
RAM[16'h721C] = 8'h00;
RAM[16'h721D] = 8'h00;
RAM[16'h721E] = 8'h00;
RAM[16'h721F] = 8'h00;
RAM[16'h7220] = 8'h00;
RAM[16'h7221] = 8'h00;
RAM[16'h7222] = 8'h00;
RAM[16'h7223] = 8'h00;
RAM[16'h7224] = 8'h00;
RAM[16'h7225] = 8'h00;
RAM[16'h7226] = 8'h00;
RAM[16'h7227] = 8'h00;
RAM[16'h7228] = 8'h00;
RAM[16'h7229] = 8'h00;
RAM[16'h722A] = 8'h00;
RAM[16'h722B] = 8'h00;
RAM[16'h722C] = 8'h00;
RAM[16'h722D] = 8'h00;
RAM[16'h722E] = 8'h00;
RAM[16'h722F] = 8'h00;
RAM[16'h7230] = 8'h00;
RAM[16'h7231] = 8'h00;
RAM[16'h7232] = 8'h00;
RAM[16'h7233] = 8'h00;
RAM[16'h7234] = 8'h00;
RAM[16'h7235] = 8'h00;
RAM[16'h7236] = 8'h00;
RAM[16'h7237] = 8'h00;
RAM[16'h7238] = 8'h00;
RAM[16'h7239] = 8'h00;
RAM[16'h723A] = 8'h00;
RAM[16'h723B] = 8'h00;
RAM[16'h723C] = 8'h00;
RAM[16'h723D] = 8'h00;
RAM[16'h723E] = 8'h00;
RAM[16'h723F] = 8'h00;
RAM[16'h7240] = 8'h00;
RAM[16'h7241] = 8'h00;
RAM[16'h7242] = 8'h00;
RAM[16'h7243] = 8'h00;
RAM[16'h7244] = 8'h00;
RAM[16'h7245] = 8'h00;
RAM[16'h7246] = 8'h00;
RAM[16'h7247] = 8'h00;
RAM[16'h7248] = 8'h00;
RAM[16'h7249] = 8'h00;
RAM[16'h724A] = 8'h00;
RAM[16'h724B] = 8'h00;
RAM[16'h724C] = 8'h00;
RAM[16'h724D] = 8'h00;
RAM[16'h724E] = 8'h00;
RAM[16'h724F] = 8'h00;
RAM[16'h7250] = 8'h00;
RAM[16'h7251] = 8'h00;
RAM[16'h7252] = 8'h00;
RAM[16'h7253] = 8'h00;
RAM[16'h7254] = 8'h00;
RAM[16'h7255] = 8'h00;
RAM[16'h7256] = 8'h00;
RAM[16'h7257] = 8'h00;
RAM[16'h7258] = 8'h00;
RAM[16'h7259] = 8'h00;
RAM[16'h725A] = 8'h00;
RAM[16'h725B] = 8'h00;
RAM[16'h725C] = 8'h00;
RAM[16'h725D] = 8'h00;
RAM[16'h725E] = 8'h00;
RAM[16'h725F] = 8'h00;
RAM[16'h7260] = 8'h00;
RAM[16'h7261] = 8'h00;
RAM[16'h7262] = 8'h00;
RAM[16'h7263] = 8'h00;
RAM[16'h7264] = 8'h00;
RAM[16'h7265] = 8'h00;
RAM[16'h7266] = 8'h00;
RAM[16'h7267] = 8'h00;
RAM[16'h7268] = 8'h00;
RAM[16'h7269] = 8'h00;
RAM[16'h726A] = 8'h00;
RAM[16'h726B] = 8'h00;
RAM[16'h726C] = 8'h00;
RAM[16'h726D] = 8'h00;
RAM[16'h726E] = 8'h00;
RAM[16'h726F] = 8'h00;
RAM[16'h7270] = 8'h00;
RAM[16'h7271] = 8'h00;
RAM[16'h7272] = 8'h00;
RAM[16'h7273] = 8'h00;
RAM[16'h7274] = 8'h00;
RAM[16'h7275] = 8'h00;
RAM[16'h7276] = 8'h00;
RAM[16'h7277] = 8'h00;
RAM[16'h7278] = 8'h00;
RAM[16'h7279] = 8'h00;
RAM[16'h727A] = 8'h00;
RAM[16'h727B] = 8'h00;
RAM[16'h727C] = 8'h00;
RAM[16'h727D] = 8'h00;
RAM[16'h727E] = 8'h00;
RAM[16'h727F] = 8'h00;
RAM[16'h7280] = 8'h00;
RAM[16'h7281] = 8'h00;
RAM[16'h7282] = 8'h00;
RAM[16'h7283] = 8'h00;
RAM[16'h7284] = 8'h00;
RAM[16'h7285] = 8'h00;
RAM[16'h7286] = 8'h00;
RAM[16'h7287] = 8'h00;
RAM[16'h7288] = 8'h00;
RAM[16'h7289] = 8'h00;
RAM[16'h728A] = 8'h00;
RAM[16'h728B] = 8'h00;
RAM[16'h728C] = 8'h00;
RAM[16'h728D] = 8'h00;
RAM[16'h728E] = 8'h00;
RAM[16'h728F] = 8'h00;
RAM[16'h7290] = 8'h00;
RAM[16'h7291] = 8'h00;
RAM[16'h7292] = 8'h00;
RAM[16'h7293] = 8'h00;
RAM[16'h7294] = 8'h00;
RAM[16'h7295] = 8'h00;
RAM[16'h7296] = 8'h00;
RAM[16'h7297] = 8'h00;
RAM[16'h7298] = 8'h00;
RAM[16'h7299] = 8'h00;
RAM[16'h729A] = 8'h00;
RAM[16'h729B] = 8'h00;
RAM[16'h729C] = 8'h00;
RAM[16'h729D] = 8'h00;
RAM[16'h729E] = 8'h00;
RAM[16'h729F] = 8'h00;
RAM[16'h72A0] = 8'h00;
RAM[16'h72A1] = 8'h00;
RAM[16'h72A2] = 8'h00;
RAM[16'h72A3] = 8'h00;
RAM[16'h72A4] = 8'h00;
RAM[16'h72A5] = 8'h00;
RAM[16'h72A6] = 8'h00;
RAM[16'h72A7] = 8'h00;
RAM[16'h72A8] = 8'h00;
RAM[16'h72A9] = 8'h00;
RAM[16'h72AA] = 8'h00;
RAM[16'h72AB] = 8'h00;
RAM[16'h72AC] = 8'h00;
RAM[16'h72AD] = 8'h00;
RAM[16'h72AE] = 8'h00;
RAM[16'h72AF] = 8'h00;
RAM[16'h72B0] = 8'h00;
RAM[16'h72B1] = 8'h00;
RAM[16'h72B2] = 8'h00;
RAM[16'h72B3] = 8'h00;
RAM[16'h72B4] = 8'h00;
RAM[16'h72B5] = 8'h00;
RAM[16'h72B6] = 8'h00;
RAM[16'h72B7] = 8'h00;
RAM[16'h72B8] = 8'h00;
RAM[16'h72B9] = 8'h00;
RAM[16'h72BA] = 8'h00;
RAM[16'h72BB] = 8'h00;
RAM[16'h72BC] = 8'h00;
RAM[16'h72BD] = 8'h00;
RAM[16'h72BE] = 8'h00;
RAM[16'h72BF] = 8'h00;
RAM[16'h72C0] = 8'h00;
RAM[16'h72C1] = 8'h00;
RAM[16'h72C2] = 8'h00;
RAM[16'h72C3] = 8'h00;
RAM[16'h72C4] = 8'h00;
RAM[16'h72C5] = 8'h00;
RAM[16'h72C6] = 8'h00;
RAM[16'h72C7] = 8'h00;
RAM[16'h72C8] = 8'h00;
RAM[16'h72C9] = 8'h00;
RAM[16'h72CA] = 8'h00;
RAM[16'h72CB] = 8'h00;
RAM[16'h72CC] = 8'h00;
RAM[16'h72CD] = 8'h00;
RAM[16'h72CE] = 8'h00;
RAM[16'h72CF] = 8'h00;
RAM[16'h72D0] = 8'h00;
RAM[16'h72D1] = 8'h00;
RAM[16'h72D2] = 8'h00;
RAM[16'h72D3] = 8'h00;
RAM[16'h72D4] = 8'h00;
RAM[16'h72D5] = 8'h00;
RAM[16'h72D6] = 8'h00;
RAM[16'h72D7] = 8'h00;
RAM[16'h72D8] = 8'h00;
RAM[16'h72D9] = 8'h00;
RAM[16'h72DA] = 8'h00;
RAM[16'h72DB] = 8'h00;
RAM[16'h72DC] = 8'h00;
RAM[16'h72DD] = 8'h00;
RAM[16'h72DE] = 8'h00;
RAM[16'h72DF] = 8'h00;
RAM[16'h72E0] = 8'h00;
RAM[16'h72E1] = 8'h00;
RAM[16'h72E2] = 8'h00;
RAM[16'h72E3] = 8'h00;
RAM[16'h72E4] = 8'h00;
RAM[16'h72E5] = 8'h00;
RAM[16'h72E6] = 8'h00;
RAM[16'h72E7] = 8'h00;
RAM[16'h72E8] = 8'h00;
RAM[16'h72E9] = 8'h00;
RAM[16'h72EA] = 8'h00;
RAM[16'h72EB] = 8'h00;
RAM[16'h72EC] = 8'h00;
RAM[16'h72ED] = 8'h00;
RAM[16'h72EE] = 8'h00;
RAM[16'h72EF] = 8'h00;
RAM[16'h72F0] = 8'h00;
RAM[16'h72F1] = 8'h00;
RAM[16'h72F2] = 8'h00;
RAM[16'h72F3] = 8'h00;
RAM[16'h72F4] = 8'h00;
RAM[16'h72F5] = 8'h00;
RAM[16'h72F6] = 8'h00;
RAM[16'h72F7] = 8'h00;
RAM[16'h72F8] = 8'h00;
RAM[16'h72F9] = 8'h00;
RAM[16'h72FA] = 8'h00;
RAM[16'h72FB] = 8'h00;
RAM[16'h72FC] = 8'h00;
RAM[16'h72FD] = 8'h00;
RAM[16'h72FE] = 8'h00;
RAM[16'h72FF] = 8'h00;
RAM[16'h7300] = 8'h00;
RAM[16'h7301] = 8'h00;
RAM[16'h7302] = 8'h00;
RAM[16'h7303] = 8'h00;
RAM[16'h7304] = 8'h00;
RAM[16'h7305] = 8'h00;
RAM[16'h7306] = 8'h00;
RAM[16'h7307] = 8'h00;
RAM[16'h7308] = 8'h00;
RAM[16'h7309] = 8'h00;
RAM[16'h730A] = 8'h00;
RAM[16'h730B] = 8'h00;
RAM[16'h730C] = 8'h00;
RAM[16'h730D] = 8'h00;
RAM[16'h730E] = 8'h00;
RAM[16'h730F] = 8'h00;
RAM[16'h7310] = 8'h00;
RAM[16'h7311] = 8'h00;
RAM[16'h7312] = 8'h00;
RAM[16'h7313] = 8'h00;
RAM[16'h7314] = 8'h00;
RAM[16'h7315] = 8'h00;
RAM[16'h7316] = 8'h00;
RAM[16'h7317] = 8'h00;
RAM[16'h7318] = 8'h00;
RAM[16'h7319] = 8'h00;
RAM[16'h731A] = 8'h00;
RAM[16'h731B] = 8'h00;
RAM[16'h731C] = 8'h00;
RAM[16'h731D] = 8'h00;
RAM[16'h731E] = 8'h00;
RAM[16'h731F] = 8'h00;
RAM[16'h7320] = 8'h00;
RAM[16'h7321] = 8'h00;
RAM[16'h7322] = 8'h00;
RAM[16'h7323] = 8'h00;
RAM[16'h7324] = 8'h00;
RAM[16'h7325] = 8'h00;
RAM[16'h7326] = 8'h00;
RAM[16'h7327] = 8'h00;
RAM[16'h7328] = 8'h00;
RAM[16'h7329] = 8'h00;
RAM[16'h732A] = 8'h00;
RAM[16'h732B] = 8'h00;
RAM[16'h732C] = 8'h00;
RAM[16'h732D] = 8'h00;
RAM[16'h732E] = 8'h00;
RAM[16'h732F] = 8'h00;
RAM[16'h7330] = 8'h00;
RAM[16'h7331] = 8'h00;
RAM[16'h7332] = 8'h00;
RAM[16'h7333] = 8'h00;
RAM[16'h7334] = 8'h00;
RAM[16'h7335] = 8'h00;
RAM[16'h7336] = 8'h00;
RAM[16'h7337] = 8'h00;
RAM[16'h7338] = 8'h00;
RAM[16'h7339] = 8'h00;
RAM[16'h733A] = 8'h00;
RAM[16'h733B] = 8'h00;
RAM[16'h733C] = 8'h00;
RAM[16'h733D] = 8'h00;
RAM[16'h733E] = 8'h00;
RAM[16'h733F] = 8'h00;
RAM[16'h7340] = 8'h00;
RAM[16'h7341] = 8'h00;
RAM[16'h7342] = 8'h00;
RAM[16'h7343] = 8'h00;
RAM[16'h7344] = 8'h00;
RAM[16'h7345] = 8'h00;
RAM[16'h7346] = 8'h00;
RAM[16'h7347] = 8'h00;
RAM[16'h7348] = 8'h00;
RAM[16'h7349] = 8'h00;
RAM[16'h734A] = 8'h00;
RAM[16'h734B] = 8'h00;
RAM[16'h734C] = 8'h00;
RAM[16'h734D] = 8'h00;
RAM[16'h734E] = 8'h00;
RAM[16'h734F] = 8'h00;
RAM[16'h7350] = 8'h00;
RAM[16'h7351] = 8'h00;
RAM[16'h7352] = 8'h00;
RAM[16'h7353] = 8'h00;
RAM[16'h7354] = 8'h00;
RAM[16'h7355] = 8'h00;
RAM[16'h7356] = 8'h00;
RAM[16'h7357] = 8'h00;
RAM[16'h7358] = 8'h00;
RAM[16'h7359] = 8'h00;
RAM[16'h735A] = 8'h00;
RAM[16'h735B] = 8'h00;
RAM[16'h735C] = 8'h00;
RAM[16'h735D] = 8'h00;
RAM[16'h735E] = 8'h00;
RAM[16'h735F] = 8'h00;
RAM[16'h7360] = 8'h00;
RAM[16'h7361] = 8'h00;
RAM[16'h7362] = 8'h00;
RAM[16'h7363] = 8'h00;
RAM[16'h7364] = 8'h00;
RAM[16'h7365] = 8'h00;
RAM[16'h7366] = 8'h00;
RAM[16'h7367] = 8'h00;
RAM[16'h7368] = 8'h00;
RAM[16'h7369] = 8'h00;
RAM[16'h736A] = 8'h00;
RAM[16'h736B] = 8'h00;
RAM[16'h736C] = 8'h00;
RAM[16'h736D] = 8'h00;
RAM[16'h736E] = 8'h00;
RAM[16'h736F] = 8'h00;
RAM[16'h7370] = 8'h00;
RAM[16'h7371] = 8'h00;
RAM[16'h7372] = 8'h00;
RAM[16'h7373] = 8'h00;
RAM[16'h7374] = 8'h00;
RAM[16'h7375] = 8'h00;
RAM[16'h7376] = 8'h00;
RAM[16'h7377] = 8'h00;
RAM[16'h7378] = 8'h00;
RAM[16'h7379] = 8'h00;
RAM[16'h737A] = 8'h00;
RAM[16'h737B] = 8'h00;
RAM[16'h737C] = 8'h00;
RAM[16'h737D] = 8'h00;
RAM[16'h737E] = 8'h00;
RAM[16'h737F] = 8'h00;
RAM[16'h7380] = 8'h00;
RAM[16'h7381] = 8'h00;
RAM[16'h7382] = 8'h00;
RAM[16'h7383] = 8'h00;
RAM[16'h7384] = 8'h00;
RAM[16'h7385] = 8'h00;
RAM[16'h7386] = 8'h00;
RAM[16'h7387] = 8'h00;
RAM[16'h7388] = 8'h00;
RAM[16'h7389] = 8'h00;
RAM[16'h738A] = 8'h00;
RAM[16'h738B] = 8'h00;
RAM[16'h738C] = 8'h00;
RAM[16'h738D] = 8'h00;
RAM[16'h738E] = 8'h00;
RAM[16'h738F] = 8'h00;
RAM[16'h7390] = 8'h00;
RAM[16'h7391] = 8'h00;
RAM[16'h7392] = 8'h00;
RAM[16'h7393] = 8'h00;
RAM[16'h7394] = 8'h00;
RAM[16'h7395] = 8'h00;
RAM[16'h7396] = 8'h00;
RAM[16'h7397] = 8'h00;
RAM[16'h7398] = 8'h00;
RAM[16'h7399] = 8'h00;
RAM[16'h739A] = 8'h00;
RAM[16'h739B] = 8'h00;
RAM[16'h739C] = 8'h00;
RAM[16'h739D] = 8'h00;
RAM[16'h739E] = 8'h00;
RAM[16'h739F] = 8'h00;
RAM[16'h73A0] = 8'h00;
RAM[16'h73A1] = 8'h00;
RAM[16'h73A2] = 8'h00;
RAM[16'h73A3] = 8'h00;
RAM[16'h73A4] = 8'h00;
RAM[16'h73A5] = 8'h00;
RAM[16'h73A6] = 8'h00;
RAM[16'h73A7] = 8'h00;
RAM[16'h73A8] = 8'h00;
RAM[16'h73A9] = 8'h00;
RAM[16'h73AA] = 8'h00;
RAM[16'h73AB] = 8'h00;
RAM[16'h73AC] = 8'h00;
RAM[16'h73AD] = 8'h00;
RAM[16'h73AE] = 8'h00;
RAM[16'h73AF] = 8'h00;
RAM[16'h73B0] = 8'h00;
RAM[16'h73B1] = 8'h00;
RAM[16'h73B2] = 8'h00;
RAM[16'h73B3] = 8'h00;
RAM[16'h73B4] = 8'h00;
RAM[16'h73B5] = 8'h00;
RAM[16'h73B6] = 8'h00;
RAM[16'h73B7] = 8'h00;
RAM[16'h73B8] = 8'h00;
RAM[16'h73B9] = 8'h00;
RAM[16'h73BA] = 8'h00;
RAM[16'h73BB] = 8'h00;
RAM[16'h73BC] = 8'h00;
RAM[16'h73BD] = 8'h00;
RAM[16'h73BE] = 8'h00;
RAM[16'h73BF] = 8'h00;
RAM[16'h73C0] = 8'h00;
RAM[16'h73C1] = 8'h00;
RAM[16'h73C2] = 8'h00;
RAM[16'h73C3] = 8'h00;
RAM[16'h73C4] = 8'h00;
RAM[16'h73C5] = 8'h00;
RAM[16'h73C6] = 8'h00;
RAM[16'h73C7] = 8'h00;
RAM[16'h73C8] = 8'h00;
RAM[16'h73C9] = 8'h00;
RAM[16'h73CA] = 8'h00;
RAM[16'h73CB] = 8'h00;
RAM[16'h73CC] = 8'h00;
RAM[16'h73CD] = 8'h00;
RAM[16'h73CE] = 8'h00;
RAM[16'h73CF] = 8'h00;
RAM[16'h73D0] = 8'h00;
RAM[16'h73D1] = 8'h00;
RAM[16'h73D2] = 8'h00;
RAM[16'h73D3] = 8'h00;
RAM[16'h73D4] = 8'h00;
RAM[16'h73D5] = 8'h00;
RAM[16'h73D6] = 8'h00;
RAM[16'h73D7] = 8'h00;
RAM[16'h73D8] = 8'h00;
RAM[16'h73D9] = 8'h00;
RAM[16'h73DA] = 8'h00;
RAM[16'h73DB] = 8'h00;
RAM[16'h73DC] = 8'h00;
RAM[16'h73DD] = 8'h00;
RAM[16'h73DE] = 8'h00;
RAM[16'h73DF] = 8'h00;
RAM[16'h73E0] = 8'h00;
RAM[16'h73E1] = 8'h00;
RAM[16'h73E2] = 8'h00;
RAM[16'h73E3] = 8'h00;
RAM[16'h73E4] = 8'h00;
RAM[16'h73E5] = 8'h00;
RAM[16'h73E6] = 8'h00;
RAM[16'h73E7] = 8'h00;
RAM[16'h73E8] = 8'h00;
RAM[16'h73E9] = 8'h00;
RAM[16'h73EA] = 8'h00;
RAM[16'h73EB] = 8'h00;
RAM[16'h73EC] = 8'h00;
RAM[16'h73ED] = 8'h00;
RAM[16'h73EE] = 8'h00;
RAM[16'h73EF] = 8'h00;
RAM[16'h73F0] = 8'h00;
RAM[16'h73F1] = 8'h00;
RAM[16'h73F2] = 8'h00;
RAM[16'h73F3] = 8'h00;
RAM[16'h73F4] = 8'h00;
RAM[16'h73F5] = 8'h00;
RAM[16'h73F6] = 8'h00;
RAM[16'h73F7] = 8'h00;
RAM[16'h73F8] = 8'h00;
RAM[16'h73F9] = 8'h00;
RAM[16'h73FA] = 8'h00;
RAM[16'h73FB] = 8'h00;
RAM[16'h73FC] = 8'h00;
RAM[16'h73FD] = 8'h00;
RAM[16'h73FE] = 8'h00;
RAM[16'h73FF] = 8'h00;
RAM[16'h7400] = 8'h00;
RAM[16'h7401] = 8'h00;
RAM[16'h7402] = 8'h00;
RAM[16'h7403] = 8'h00;
RAM[16'h7404] = 8'h00;
RAM[16'h7405] = 8'h00;
RAM[16'h7406] = 8'h00;
RAM[16'h7407] = 8'h00;
RAM[16'h7408] = 8'h00;
RAM[16'h7409] = 8'h00;
RAM[16'h740A] = 8'h00;
RAM[16'h740B] = 8'h00;
RAM[16'h740C] = 8'h00;
RAM[16'h740D] = 8'h00;
RAM[16'h740E] = 8'h00;
RAM[16'h740F] = 8'h00;
RAM[16'h7410] = 8'h00;
RAM[16'h7411] = 8'h00;
RAM[16'h7412] = 8'h00;
RAM[16'h7413] = 8'h00;
RAM[16'h7414] = 8'h00;
RAM[16'h7415] = 8'h00;
RAM[16'h7416] = 8'h00;
RAM[16'h7417] = 8'h00;
RAM[16'h7418] = 8'h00;
RAM[16'h7419] = 8'h00;
RAM[16'h741A] = 8'h00;
RAM[16'h741B] = 8'h00;
RAM[16'h741C] = 8'h00;
RAM[16'h741D] = 8'h00;
RAM[16'h741E] = 8'h00;
RAM[16'h741F] = 8'h00;
RAM[16'h7420] = 8'h00;
RAM[16'h7421] = 8'h00;
RAM[16'h7422] = 8'h00;
RAM[16'h7423] = 8'h00;
RAM[16'h7424] = 8'h00;
RAM[16'h7425] = 8'h00;
RAM[16'h7426] = 8'h00;
RAM[16'h7427] = 8'h00;
RAM[16'h7428] = 8'h00;
RAM[16'h7429] = 8'h00;
RAM[16'h742A] = 8'h00;
RAM[16'h742B] = 8'h00;
RAM[16'h742C] = 8'h00;
RAM[16'h742D] = 8'h00;
RAM[16'h742E] = 8'h00;
RAM[16'h742F] = 8'h00;
RAM[16'h7430] = 8'h00;
RAM[16'h7431] = 8'h00;
RAM[16'h7432] = 8'h00;
RAM[16'h7433] = 8'h00;
RAM[16'h7434] = 8'h00;
RAM[16'h7435] = 8'h00;
RAM[16'h7436] = 8'h00;
RAM[16'h7437] = 8'h00;
RAM[16'h7438] = 8'h00;
RAM[16'h7439] = 8'h00;
RAM[16'h743A] = 8'h00;
RAM[16'h743B] = 8'h00;
RAM[16'h743C] = 8'h00;
RAM[16'h743D] = 8'h00;
RAM[16'h743E] = 8'h00;
RAM[16'h743F] = 8'h00;
RAM[16'h7440] = 8'h00;
RAM[16'h7441] = 8'h00;
RAM[16'h7442] = 8'h00;
RAM[16'h7443] = 8'h00;
RAM[16'h7444] = 8'h00;
RAM[16'h7445] = 8'h00;
RAM[16'h7446] = 8'h00;
RAM[16'h7447] = 8'h00;
RAM[16'h7448] = 8'h00;
RAM[16'h7449] = 8'h00;
RAM[16'h744A] = 8'h00;
RAM[16'h744B] = 8'h00;
RAM[16'h744C] = 8'h00;
RAM[16'h744D] = 8'h00;
RAM[16'h744E] = 8'h00;
RAM[16'h744F] = 8'h00;
RAM[16'h7450] = 8'h00;
RAM[16'h7451] = 8'h00;
RAM[16'h7452] = 8'h00;
RAM[16'h7453] = 8'h00;
RAM[16'h7454] = 8'h00;
RAM[16'h7455] = 8'h00;
RAM[16'h7456] = 8'h00;
RAM[16'h7457] = 8'h00;
RAM[16'h7458] = 8'h00;
RAM[16'h7459] = 8'h00;
RAM[16'h745A] = 8'h00;
RAM[16'h745B] = 8'h00;
RAM[16'h745C] = 8'h00;
RAM[16'h745D] = 8'h00;
RAM[16'h745E] = 8'h00;
RAM[16'h745F] = 8'h00;
RAM[16'h7460] = 8'h00;
RAM[16'h7461] = 8'h00;
RAM[16'h7462] = 8'h00;
RAM[16'h7463] = 8'h00;
RAM[16'h7464] = 8'h00;
RAM[16'h7465] = 8'h00;
RAM[16'h7466] = 8'h00;
RAM[16'h7467] = 8'h00;
RAM[16'h7468] = 8'h00;
RAM[16'h7469] = 8'h00;
RAM[16'h746A] = 8'h00;
RAM[16'h746B] = 8'h00;
RAM[16'h746C] = 8'h00;
RAM[16'h746D] = 8'h00;
RAM[16'h746E] = 8'h00;
RAM[16'h746F] = 8'h00;
RAM[16'h7470] = 8'h00;
RAM[16'h7471] = 8'h00;
RAM[16'h7472] = 8'h00;
RAM[16'h7473] = 8'h00;
RAM[16'h7474] = 8'h00;
RAM[16'h7475] = 8'h00;
RAM[16'h7476] = 8'h00;
RAM[16'h7477] = 8'h00;
RAM[16'h7478] = 8'h00;
RAM[16'h7479] = 8'h00;
RAM[16'h747A] = 8'h00;
RAM[16'h747B] = 8'h00;
RAM[16'h747C] = 8'h00;
RAM[16'h747D] = 8'h00;
RAM[16'h747E] = 8'h00;
RAM[16'h747F] = 8'h00;
RAM[16'h7480] = 8'h00;
RAM[16'h7481] = 8'h00;
RAM[16'h7482] = 8'h00;
RAM[16'h7483] = 8'h00;
RAM[16'h7484] = 8'h00;
RAM[16'h7485] = 8'h00;
RAM[16'h7486] = 8'h00;
RAM[16'h7487] = 8'h00;
RAM[16'h7488] = 8'h00;
RAM[16'h7489] = 8'h00;
RAM[16'h748A] = 8'h00;
RAM[16'h748B] = 8'h00;
RAM[16'h748C] = 8'h00;
RAM[16'h748D] = 8'h00;
RAM[16'h748E] = 8'h00;
RAM[16'h748F] = 8'h00;
RAM[16'h7490] = 8'h00;
RAM[16'h7491] = 8'h00;
RAM[16'h7492] = 8'h00;
RAM[16'h7493] = 8'h00;
RAM[16'h7494] = 8'h00;
RAM[16'h7495] = 8'h00;
RAM[16'h7496] = 8'h00;
RAM[16'h7497] = 8'h00;
RAM[16'h7498] = 8'h00;
RAM[16'h7499] = 8'h00;
RAM[16'h749A] = 8'h00;
RAM[16'h749B] = 8'h00;
RAM[16'h749C] = 8'h00;
RAM[16'h749D] = 8'h00;
RAM[16'h749E] = 8'h00;
RAM[16'h749F] = 8'h00;
RAM[16'h74A0] = 8'h00;
RAM[16'h74A1] = 8'h00;
RAM[16'h74A2] = 8'h00;
RAM[16'h74A3] = 8'h00;
RAM[16'h74A4] = 8'h00;
RAM[16'h74A5] = 8'h00;
RAM[16'h74A6] = 8'h00;
RAM[16'h74A7] = 8'h00;
RAM[16'h74A8] = 8'h00;
RAM[16'h74A9] = 8'h00;
RAM[16'h74AA] = 8'h00;
RAM[16'h74AB] = 8'h00;
RAM[16'h74AC] = 8'h00;
RAM[16'h74AD] = 8'h00;
RAM[16'h74AE] = 8'h00;
RAM[16'h74AF] = 8'h00;
RAM[16'h74B0] = 8'h00;
RAM[16'h74B1] = 8'h00;
RAM[16'h74B2] = 8'h00;
RAM[16'h74B3] = 8'h00;
RAM[16'h74B4] = 8'h00;
RAM[16'h74B5] = 8'h00;
RAM[16'h74B6] = 8'h00;
RAM[16'h74B7] = 8'h00;
RAM[16'h74B8] = 8'h00;
RAM[16'h74B9] = 8'h00;
RAM[16'h74BA] = 8'h00;
RAM[16'h74BB] = 8'h00;
RAM[16'h74BC] = 8'h00;
RAM[16'h74BD] = 8'h00;
RAM[16'h74BE] = 8'h00;
RAM[16'h74BF] = 8'h00;
RAM[16'h74C0] = 8'h00;
RAM[16'h74C1] = 8'h00;
RAM[16'h74C2] = 8'h00;
RAM[16'h74C3] = 8'h00;
RAM[16'h74C4] = 8'h00;
RAM[16'h74C5] = 8'h00;
RAM[16'h74C6] = 8'h00;
RAM[16'h74C7] = 8'h00;
RAM[16'h74C8] = 8'h00;
RAM[16'h74C9] = 8'h00;
RAM[16'h74CA] = 8'h00;
RAM[16'h74CB] = 8'h00;
RAM[16'h74CC] = 8'h00;
RAM[16'h74CD] = 8'h00;
RAM[16'h74CE] = 8'h00;
RAM[16'h74CF] = 8'h00;
RAM[16'h74D0] = 8'h00;
RAM[16'h74D1] = 8'h00;
RAM[16'h74D2] = 8'h00;
RAM[16'h74D3] = 8'h00;
RAM[16'h74D4] = 8'h00;
RAM[16'h74D5] = 8'h00;
RAM[16'h74D6] = 8'h00;
RAM[16'h74D7] = 8'h00;
RAM[16'h74D8] = 8'h00;
RAM[16'h74D9] = 8'h00;
RAM[16'h74DA] = 8'h00;
RAM[16'h74DB] = 8'h00;
RAM[16'h74DC] = 8'h00;
RAM[16'h74DD] = 8'h00;
RAM[16'h74DE] = 8'h00;
RAM[16'h74DF] = 8'h00;
RAM[16'h74E0] = 8'h00;
RAM[16'h74E1] = 8'h00;
RAM[16'h74E2] = 8'h00;
RAM[16'h74E3] = 8'h00;
RAM[16'h74E4] = 8'h00;
RAM[16'h74E5] = 8'h00;
RAM[16'h74E6] = 8'h00;
RAM[16'h74E7] = 8'h00;
RAM[16'h74E8] = 8'h00;
RAM[16'h74E9] = 8'h00;
RAM[16'h74EA] = 8'h00;
RAM[16'h74EB] = 8'h00;
RAM[16'h74EC] = 8'h00;
RAM[16'h74ED] = 8'h00;
RAM[16'h74EE] = 8'h00;
RAM[16'h74EF] = 8'h00;
RAM[16'h74F0] = 8'h00;
RAM[16'h74F1] = 8'h00;
RAM[16'h74F2] = 8'h00;
RAM[16'h74F3] = 8'h00;
RAM[16'h74F4] = 8'h00;
RAM[16'h74F5] = 8'h00;
RAM[16'h74F6] = 8'h00;
RAM[16'h74F7] = 8'h00;
RAM[16'h74F8] = 8'h00;
RAM[16'h74F9] = 8'h00;
RAM[16'h74FA] = 8'h00;
RAM[16'h74FB] = 8'h00;
RAM[16'h74FC] = 8'h00;
RAM[16'h74FD] = 8'h00;
RAM[16'h74FE] = 8'h00;
RAM[16'h74FF] = 8'h00;
RAM[16'h7500] = 8'h00;
RAM[16'h7501] = 8'h00;
RAM[16'h7502] = 8'h00;
RAM[16'h7503] = 8'h00;
RAM[16'h7504] = 8'h00;
RAM[16'h7505] = 8'h00;
RAM[16'h7506] = 8'h00;
RAM[16'h7507] = 8'h00;
RAM[16'h7508] = 8'h00;
RAM[16'h7509] = 8'h00;
RAM[16'h750A] = 8'h00;
RAM[16'h750B] = 8'h00;
RAM[16'h750C] = 8'h00;
RAM[16'h750D] = 8'h00;
RAM[16'h750E] = 8'h00;
RAM[16'h750F] = 8'h00;
RAM[16'h7510] = 8'h00;
RAM[16'h7511] = 8'h00;
RAM[16'h7512] = 8'h00;
RAM[16'h7513] = 8'h00;
RAM[16'h7514] = 8'h00;
RAM[16'h7515] = 8'h00;
RAM[16'h7516] = 8'h00;
RAM[16'h7517] = 8'h00;
RAM[16'h7518] = 8'h00;
RAM[16'h7519] = 8'h00;
RAM[16'h751A] = 8'h00;
RAM[16'h751B] = 8'h00;
RAM[16'h751C] = 8'h00;
RAM[16'h751D] = 8'h00;
RAM[16'h751E] = 8'h00;
RAM[16'h751F] = 8'h00;
RAM[16'h7520] = 8'h00;
RAM[16'h7521] = 8'h00;
RAM[16'h7522] = 8'h00;
RAM[16'h7523] = 8'h00;
RAM[16'h7524] = 8'h00;
RAM[16'h7525] = 8'h00;
RAM[16'h7526] = 8'h00;
RAM[16'h7527] = 8'h00;
RAM[16'h7528] = 8'h00;
RAM[16'h7529] = 8'h00;
RAM[16'h752A] = 8'h00;
RAM[16'h752B] = 8'h00;
RAM[16'h752C] = 8'h00;
RAM[16'h752D] = 8'h00;
RAM[16'h752E] = 8'h00;
RAM[16'h752F] = 8'h00;
RAM[16'h7530] = 8'h00;
RAM[16'h7531] = 8'h00;
RAM[16'h7532] = 8'h00;
RAM[16'h7533] = 8'h00;
RAM[16'h7534] = 8'h00;
RAM[16'h7535] = 8'h00;
RAM[16'h7536] = 8'h00;
RAM[16'h7537] = 8'h00;
RAM[16'h7538] = 8'h00;
RAM[16'h7539] = 8'h00;
RAM[16'h753A] = 8'h00;
RAM[16'h753B] = 8'h00;
RAM[16'h753C] = 8'h00;
RAM[16'h753D] = 8'h00;
RAM[16'h753E] = 8'h00;
RAM[16'h753F] = 8'h00;
RAM[16'h7540] = 8'h00;
RAM[16'h7541] = 8'h00;
RAM[16'h7542] = 8'h00;
RAM[16'h7543] = 8'h00;
RAM[16'h7544] = 8'h00;
RAM[16'h7545] = 8'h00;
RAM[16'h7546] = 8'h00;
RAM[16'h7547] = 8'h00;
RAM[16'h7548] = 8'h00;
RAM[16'h7549] = 8'h00;
RAM[16'h754A] = 8'h00;
RAM[16'h754B] = 8'h00;
RAM[16'h754C] = 8'h00;
RAM[16'h754D] = 8'h00;
RAM[16'h754E] = 8'h00;
RAM[16'h754F] = 8'h00;
RAM[16'h7550] = 8'h00;
RAM[16'h7551] = 8'h00;
RAM[16'h7552] = 8'h00;
RAM[16'h7553] = 8'h00;
RAM[16'h7554] = 8'h00;
RAM[16'h7555] = 8'h00;
RAM[16'h7556] = 8'h00;
RAM[16'h7557] = 8'h00;
RAM[16'h7558] = 8'h00;
RAM[16'h7559] = 8'h00;
RAM[16'h755A] = 8'h00;
RAM[16'h755B] = 8'h00;
RAM[16'h755C] = 8'h00;
RAM[16'h755D] = 8'h00;
RAM[16'h755E] = 8'h00;
RAM[16'h755F] = 8'h00;
RAM[16'h7560] = 8'h00;
RAM[16'h7561] = 8'h00;
RAM[16'h7562] = 8'h00;
RAM[16'h7563] = 8'h00;
RAM[16'h7564] = 8'h00;
RAM[16'h7565] = 8'h00;
RAM[16'h7566] = 8'h00;
RAM[16'h7567] = 8'h00;
RAM[16'h7568] = 8'h00;
RAM[16'h7569] = 8'h00;
RAM[16'h756A] = 8'h00;
RAM[16'h756B] = 8'h00;
RAM[16'h756C] = 8'h00;
RAM[16'h756D] = 8'h00;
RAM[16'h756E] = 8'h00;
RAM[16'h756F] = 8'h00;
RAM[16'h7570] = 8'h00;
RAM[16'h7571] = 8'h00;
RAM[16'h7572] = 8'h00;
RAM[16'h7573] = 8'h00;
RAM[16'h7574] = 8'h00;
RAM[16'h7575] = 8'h00;
RAM[16'h7576] = 8'h00;
RAM[16'h7577] = 8'h00;
RAM[16'h7578] = 8'h00;
RAM[16'h7579] = 8'h00;
RAM[16'h757A] = 8'h00;
RAM[16'h757B] = 8'h00;
RAM[16'h757C] = 8'h00;
RAM[16'h757D] = 8'h00;
RAM[16'h757E] = 8'h00;
RAM[16'h757F] = 8'h00;
RAM[16'h7580] = 8'h00;
RAM[16'h7581] = 8'h00;
RAM[16'h7582] = 8'h00;
RAM[16'h7583] = 8'h00;
RAM[16'h7584] = 8'h00;
RAM[16'h7585] = 8'h00;
RAM[16'h7586] = 8'h00;
RAM[16'h7587] = 8'h00;
RAM[16'h7588] = 8'h00;
RAM[16'h7589] = 8'h00;
RAM[16'h758A] = 8'h00;
RAM[16'h758B] = 8'h00;
RAM[16'h758C] = 8'h00;
RAM[16'h758D] = 8'h00;
RAM[16'h758E] = 8'h00;
RAM[16'h758F] = 8'h00;
RAM[16'h7590] = 8'h00;
RAM[16'h7591] = 8'h00;
RAM[16'h7592] = 8'h00;
RAM[16'h7593] = 8'h00;
RAM[16'h7594] = 8'h00;
RAM[16'h7595] = 8'h00;
RAM[16'h7596] = 8'h00;
RAM[16'h7597] = 8'h00;
RAM[16'h7598] = 8'h00;
RAM[16'h7599] = 8'h00;
RAM[16'h759A] = 8'h00;
RAM[16'h759B] = 8'h00;
RAM[16'h759C] = 8'h00;
RAM[16'h759D] = 8'h00;
RAM[16'h759E] = 8'h00;
RAM[16'h759F] = 8'h00;
RAM[16'h75A0] = 8'h00;
RAM[16'h75A1] = 8'h00;
RAM[16'h75A2] = 8'h00;
RAM[16'h75A3] = 8'h00;
RAM[16'h75A4] = 8'h00;
RAM[16'h75A5] = 8'h00;
RAM[16'h75A6] = 8'h00;
RAM[16'h75A7] = 8'h00;
RAM[16'h75A8] = 8'h00;
RAM[16'h75A9] = 8'h00;
RAM[16'h75AA] = 8'h00;
RAM[16'h75AB] = 8'h00;
RAM[16'h75AC] = 8'h00;
RAM[16'h75AD] = 8'h00;
RAM[16'h75AE] = 8'h00;
RAM[16'h75AF] = 8'h00;
RAM[16'h75B0] = 8'h00;
RAM[16'h75B1] = 8'h00;
RAM[16'h75B2] = 8'h00;
RAM[16'h75B3] = 8'h00;
RAM[16'h75B4] = 8'h00;
RAM[16'h75B5] = 8'h00;
RAM[16'h75B6] = 8'h00;
RAM[16'h75B7] = 8'h00;
RAM[16'h75B8] = 8'h00;
RAM[16'h75B9] = 8'h00;
RAM[16'h75BA] = 8'h00;
RAM[16'h75BB] = 8'h00;
RAM[16'h75BC] = 8'h00;
RAM[16'h75BD] = 8'h00;
RAM[16'h75BE] = 8'h00;
RAM[16'h75BF] = 8'h00;
RAM[16'h75C0] = 8'h00;
RAM[16'h75C1] = 8'h00;
RAM[16'h75C2] = 8'h00;
RAM[16'h75C3] = 8'h00;
RAM[16'h75C4] = 8'h00;
RAM[16'h75C5] = 8'h00;
RAM[16'h75C6] = 8'h00;
RAM[16'h75C7] = 8'h00;
RAM[16'h75C8] = 8'h00;
RAM[16'h75C9] = 8'h00;
RAM[16'h75CA] = 8'h00;
RAM[16'h75CB] = 8'h00;
RAM[16'h75CC] = 8'h00;
RAM[16'h75CD] = 8'h00;
RAM[16'h75CE] = 8'h00;
RAM[16'h75CF] = 8'h00;
RAM[16'h75D0] = 8'h00;
RAM[16'h75D1] = 8'h00;
RAM[16'h75D2] = 8'h00;
RAM[16'h75D3] = 8'h00;
RAM[16'h75D4] = 8'h00;
RAM[16'h75D5] = 8'h00;
RAM[16'h75D6] = 8'h00;
RAM[16'h75D7] = 8'h00;
RAM[16'h75D8] = 8'h00;
RAM[16'h75D9] = 8'h00;
RAM[16'h75DA] = 8'h00;
RAM[16'h75DB] = 8'h00;
RAM[16'h75DC] = 8'h00;
RAM[16'h75DD] = 8'h00;
RAM[16'h75DE] = 8'h00;
RAM[16'h75DF] = 8'h00;
RAM[16'h75E0] = 8'h00;
RAM[16'h75E1] = 8'h00;
RAM[16'h75E2] = 8'h00;
RAM[16'h75E3] = 8'h00;
RAM[16'h75E4] = 8'h00;
RAM[16'h75E5] = 8'h00;
RAM[16'h75E6] = 8'h00;
RAM[16'h75E7] = 8'h00;
RAM[16'h75E8] = 8'h00;
RAM[16'h75E9] = 8'h00;
RAM[16'h75EA] = 8'h00;
RAM[16'h75EB] = 8'h00;
RAM[16'h75EC] = 8'h00;
RAM[16'h75ED] = 8'h00;
RAM[16'h75EE] = 8'h00;
RAM[16'h75EF] = 8'h00;
RAM[16'h75F0] = 8'h00;
RAM[16'h75F1] = 8'h00;
RAM[16'h75F2] = 8'h00;
RAM[16'h75F3] = 8'h00;
RAM[16'h75F4] = 8'h00;
RAM[16'h75F5] = 8'h00;
RAM[16'h75F6] = 8'h00;
RAM[16'h75F7] = 8'h00;
RAM[16'h75F8] = 8'h00;
RAM[16'h75F9] = 8'h00;
RAM[16'h75FA] = 8'h00;
RAM[16'h75FB] = 8'h00;
RAM[16'h75FC] = 8'h00;
RAM[16'h75FD] = 8'h00;
RAM[16'h75FE] = 8'h00;
RAM[16'h75FF] = 8'h00;
RAM[16'h7600] = 8'h00;
RAM[16'h7601] = 8'h00;
RAM[16'h7602] = 8'h00;
RAM[16'h7603] = 8'h00;
RAM[16'h7604] = 8'h00;
RAM[16'h7605] = 8'h00;
RAM[16'h7606] = 8'h00;
RAM[16'h7607] = 8'h00;
RAM[16'h7608] = 8'h00;
RAM[16'h7609] = 8'h00;
RAM[16'h760A] = 8'h00;
RAM[16'h760B] = 8'h00;
RAM[16'h760C] = 8'h00;
RAM[16'h760D] = 8'h00;
RAM[16'h760E] = 8'h00;
RAM[16'h760F] = 8'h00;
RAM[16'h7610] = 8'h00;
RAM[16'h7611] = 8'h00;
RAM[16'h7612] = 8'h00;
RAM[16'h7613] = 8'h00;
RAM[16'h7614] = 8'h00;
RAM[16'h7615] = 8'h00;
RAM[16'h7616] = 8'h00;
RAM[16'h7617] = 8'h00;
RAM[16'h7618] = 8'h00;
RAM[16'h7619] = 8'h00;
RAM[16'h761A] = 8'h00;
RAM[16'h761B] = 8'h00;
RAM[16'h761C] = 8'h00;
RAM[16'h761D] = 8'h00;
RAM[16'h761E] = 8'h00;
RAM[16'h761F] = 8'h00;
RAM[16'h7620] = 8'h00;
RAM[16'h7621] = 8'h00;
RAM[16'h7622] = 8'h00;
RAM[16'h7623] = 8'h00;
RAM[16'h7624] = 8'h00;
RAM[16'h7625] = 8'h00;
RAM[16'h7626] = 8'h00;
RAM[16'h7627] = 8'h00;
RAM[16'h7628] = 8'h00;
RAM[16'h7629] = 8'h00;
RAM[16'h762A] = 8'h00;
RAM[16'h762B] = 8'h00;
RAM[16'h762C] = 8'h00;
RAM[16'h762D] = 8'h00;
RAM[16'h762E] = 8'h00;
RAM[16'h762F] = 8'h00;
RAM[16'h7630] = 8'h00;
RAM[16'h7631] = 8'h00;
RAM[16'h7632] = 8'h00;
RAM[16'h7633] = 8'h00;
RAM[16'h7634] = 8'h00;
RAM[16'h7635] = 8'h00;
RAM[16'h7636] = 8'h00;
RAM[16'h7637] = 8'h00;
RAM[16'h7638] = 8'h00;
RAM[16'h7639] = 8'h00;
RAM[16'h763A] = 8'h00;
RAM[16'h763B] = 8'h00;
RAM[16'h763C] = 8'h00;
RAM[16'h763D] = 8'h00;
RAM[16'h763E] = 8'h00;
RAM[16'h763F] = 8'h00;
RAM[16'h7640] = 8'h00;
RAM[16'h7641] = 8'h00;
RAM[16'h7642] = 8'h00;
RAM[16'h7643] = 8'h00;
RAM[16'h7644] = 8'h00;
RAM[16'h7645] = 8'h00;
RAM[16'h7646] = 8'h00;
RAM[16'h7647] = 8'h00;
RAM[16'h7648] = 8'h00;
RAM[16'h7649] = 8'h00;
RAM[16'h764A] = 8'h00;
RAM[16'h764B] = 8'h00;
RAM[16'h764C] = 8'h00;
RAM[16'h764D] = 8'h00;
RAM[16'h764E] = 8'h00;
RAM[16'h764F] = 8'h00;
RAM[16'h7650] = 8'h00;
RAM[16'h7651] = 8'h00;
RAM[16'h7652] = 8'h00;
RAM[16'h7653] = 8'h00;
RAM[16'h7654] = 8'h00;
RAM[16'h7655] = 8'h00;
RAM[16'h7656] = 8'h00;
RAM[16'h7657] = 8'h00;
RAM[16'h7658] = 8'h00;
RAM[16'h7659] = 8'h00;
RAM[16'h765A] = 8'h00;
RAM[16'h765B] = 8'h00;
RAM[16'h765C] = 8'h00;
RAM[16'h765D] = 8'h00;
RAM[16'h765E] = 8'h00;
RAM[16'h765F] = 8'h00;
RAM[16'h7660] = 8'h00;
RAM[16'h7661] = 8'h00;
RAM[16'h7662] = 8'h00;
RAM[16'h7663] = 8'h00;
RAM[16'h7664] = 8'h00;
RAM[16'h7665] = 8'h00;
RAM[16'h7666] = 8'h00;
RAM[16'h7667] = 8'h00;
RAM[16'h7668] = 8'h00;
RAM[16'h7669] = 8'h00;
RAM[16'h766A] = 8'h00;
RAM[16'h766B] = 8'h00;
RAM[16'h766C] = 8'h00;
RAM[16'h766D] = 8'h00;
RAM[16'h766E] = 8'h00;
RAM[16'h766F] = 8'h00;
RAM[16'h7670] = 8'h00;
RAM[16'h7671] = 8'h00;
RAM[16'h7672] = 8'h00;
RAM[16'h7673] = 8'h00;
RAM[16'h7674] = 8'h00;
RAM[16'h7675] = 8'h00;
RAM[16'h7676] = 8'h00;
RAM[16'h7677] = 8'h00;
RAM[16'h7678] = 8'h00;
RAM[16'h7679] = 8'h00;
RAM[16'h767A] = 8'h00;
RAM[16'h767B] = 8'h00;
RAM[16'h767C] = 8'h00;
RAM[16'h767D] = 8'h00;
RAM[16'h767E] = 8'h00;
RAM[16'h767F] = 8'h00;
RAM[16'h7680] = 8'h00;
RAM[16'h7681] = 8'h00;
RAM[16'h7682] = 8'h00;
RAM[16'h7683] = 8'h00;
RAM[16'h7684] = 8'h00;
RAM[16'h7685] = 8'h00;
RAM[16'h7686] = 8'h00;
RAM[16'h7687] = 8'h00;
RAM[16'h7688] = 8'h00;
RAM[16'h7689] = 8'h00;
RAM[16'h768A] = 8'h00;
RAM[16'h768B] = 8'h00;
RAM[16'h768C] = 8'h00;
RAM[16'h768D] = 8'h00;
RAM[16'h768E] = 8'h00;
RAM[16'h768F] = 8'h00;
RAM[16'h7690] = 8'h00;
RAM[16'h7691] = 8'h00;
RAM[16'h7692] = 8'h00;
RAM[16'h7693] = 8'h00;
RAM[16'h7694] = 8'h00;
RAM[16'h7695] = 8'h00;
RAM[16'h7696] = 8'h00;
RAM[16'h7697] = 8'h00;
RAM[16'h7698] = 8'h00;
RAM[16'h7699] = 8'h00;
RAM[16'h769A] = 8'h00;
RAM[16'h769B] = 8'h00;
RAM[16'h769C] = 8'h00;
RAM[16'h769D] = 8'h00;
RAM[16'h769E] = 8'h00;
RAM[16'h769F] = 8'h00;
RAM[16'h76A0] = 8'h00;
RAM[16'h76A1] = 8'h00;
RAM[16'h76A2] = 8'h00;
RAM[16'h76A3] = 8'h00;
RAM[16'h76A4] = 8'h00;
RAM[16'h76A5] = 8'h00;
RAM[16'h76A6] = 8'h00;
RAM[16'h76A7] = 8'h00;
RAM[16'h76A8] = 8'h00;
RAM[16'h76A9] = 8'h00;
RAM[16'h76AA] = 8'h00;
RAM[16'h76AB] = 8'h00;
RAM[16'h76AC] = 8'h00;
RAM[16'h76AD] = 8'h00;
RAM[16'h76AE] = 8'h00;
RAM[16'h76AF] = 8'h00;
RAM[16'h76B0] = 8'h00;
RAM[16'h76B1] = 8'h00;
RAM[16'h76B2] = 8'h00;
RAM[16'h76B3] = 8'h00;
RAM[16'h76B4] = 8'h00;
RAM[16'h76B5] = 8'h00;
RAM[16'h76B6] = 8'h00;
RAM[16'h76B7] = 8'h00;
RAM[16'h76B8] = 8'h00;
RAM[16'h76B9] = 8'h00;
RAM[16'h76BA] = 8'h00;
RAM[16'h76BB] = 8'h00;
RAM[16'h76BC] = 8'h00;
RAM[16'h76BD] = 8'h00;
RAM[16'h76BE] = 8'h00;
RAM[16'h76BF] = 8'h00;
RAM[16'h76C0] = 8'h00;
RAM[16'h76C1] = 8'h00;
RAM[16'h76C2] = 8'h00;
RAM[16'h76C3] = 8'h00;
RAM[16'h76C4] = 8'h00;
RAM[16'h76C5] = 8'h00;
RAM[16'h76C6] = 8'h00;
RAM[16'h76C7] = 8'h00;
RAM[16'h76C8] = 8'h00;
RAM[16'h76C9] = 8'h00;
RAM[16'h76CA] = 8'h00;
RAM[16'h76CB] = 8'h00;
RAM[16'h76CC] = 8'h00;
RAM[16'h76CD] = 8'h00;
RAM[16'h76CE] = 8'h00;
RAM[16'h76CF] = 8'h00;
RAM[16'h76D0] = 8'h00;
RAM[16'h76D1] = 8'h00;
RAM[16'h76D2] = 8'h00;
RAM[16'h76D3] = 8'h00;
RAM[16'h76D4] = 8'h00;
RAM[16'h76D5] = 8'h00;
RAM[16'h76D6] = 8'h00;
RAM[16'h76D7] = 8'h00;
RAM[16'h76D8] = 8'h00;
RAM[16'h76D9] = 8'h00;
RAM[16'h76DA] = 8'h00;
RAM[16'h76DB] = 8'h00;
RAM[16'h76DC] = 8'h00;
RAM[16'h76DD] = 8'h00;
RAM[16'h76DE] = 8'h00;
RAM[16'h76DF] = 8'h00;
RAM[16'h76E0] = 8'h00;
RAM[16'h76E1] = 8'h00;
RAM[16'h76E2] = 8'h00;
RAM[16'h76E3] = 8'h00;
RAM[16'h76E4] = 8'h00;
RAM[16'h76E5] = 8'h00;
RAM[16'h76E6] = 8'h00;
RAM[16'h76E7] = 8'h00;
RAM[16'h76E8] = 8'h00;
RAM[16'h76E9] = 8'h00;
RAM[16'h76EA] = 8'h00;
RAM[16'h76EB] = 8'h00;
RAM[16'h76EC] = 8'h00;
RAM[16'h76ED] = 8'h00;
RAM[16'h76EE] = 8'h00;
RAM[16'h76EF] = 8'h00;
RAM[16'h76F0] = 8'h00;
RAM[16'h76F1] = 8'h00;
RAM[16'h76F2] = 8'h00;
RAM[16'h76F3] = 8'h00;
RAM[16'h76F4] = 8'h00;
RAM[16'h76F5] = 8'h00;
RAM[16'h76F6] = 8'h00;
RAM[16'h76F7] = 8'h00;
RAM[16'h76F8] = 8'h00;
RAM[16'h76F9] = 8'h00;
RAM[16'h76FA] = 8'h00;
RAM[16'h76FB] = 8'h00;
RAM[16'h76FC] = 8'h00;
RAM[16'h76FD] = 8'h00;
RAM[16'h76FE] = 8'h00;
RAM[16'h76FF] = 8'h00;
RAM[16'h7700] = 8'h00;
RAM[16'h7701] = 8'h00;
RAM[16'h7702] = 8'h00;
RAM[16'h7703] = 8'h00;
RAM[16'h7704] = 8'h00;
RAM[16'h7705] = 8'h00;
RAM[16'h7706] = 8'h00;
RAM[16'h7707] = 8'h00;
RAM[16'h7708] = 8'h00;
RAM[16'h7709] = 8'h00;
RAM[16'h770A] = 8'h00;
RAM[16'h770B] = 8'h00;
RAM[16'h770C] = 8'h00;
RAM[16'h770D] = 8'h00;
RAM[16'h770E] = 8'h00;
RAM[16'h770F] = 8'h00;
RAM[16'h7710] = 8'h00;
RAM[16'h7711] = 8'h00;
RAM[16'h7712] = 8'h00;
RAM[16'h7713] = 8'h00;
RAM[16'h7714] = 8'h00;
RAM[16'h7715] = 8'h00;
RAM[16'h7716] = 8'h00;
RAM[16'h7717] = 8'h00;
RAM[16'h7718] = 8'h00;
RAM[16'h7719] = 8'h00;
RAM[16'h771A] = 8'h00;
RAM[16'h771B] = 8'h00;
RAM[16'h771C] = 8'h00;
RAM[16'h771D] = 8'h00;
RAM[16'h771E] = 8'h00;
RAM[16'h771F] = 8'h00;
RAM[16'h7720] = 8'h00;
RAM[16'h7721] = 8'h00;
RAM[16'h7722] = 8'h00;
RAM[16'h7723] = 8'h00;
RAM[16'h7724] = 8'h00;
RAM[16'h7725] = 8'h00;
RAM[16'h7726] = 8'h00;
RAM[16'h7727] = 8'h00;
RAM[16'h7728] = 8'h00;
RAM[16'h7729] = 8'h00;
RAM[16'h772A] = 8'h00;
RAM[16'h772B] = 8'h00;
RAM[16'h772C] = 8'h00;
RAM[16'h772D] = 8'h00;
RAM[16'h772E] = 8'h00;
RAM[16'h772F] = 8'h00;
RAM[16'h7730] = 8'h00;
RAM[16'h7731] = 8'h00;
RAM[16'h7732] = 8'h00;
RAM[16'h7733] = 8'h00;
RAM[16'h7734] = 8'h00;
RAM[16'h7735] = 8'h00;
RAM[16'h7736] = 8'h00;
RAM[16'h7737] = 8'h00;
RAM[16'h7738] = 8'h00;
RAM[16'h7739] = 8'h00;
RAM[16'h773A] = 8'h00;
RAM[16'h773B] = 8'h00;
RAM[16'h773C] = 8'h00;
RAM[16'h773D] = 8'h00;
RAM[16'h773E] = 8'h00;
RAM[16'h773F] = 8'h00;
RAM[16'h7740] = 8'h00;
RAM[16'h7741] = 8'h00;
RAM[16'h7742] = 8'h00;
RAM[16'h7743] = 8'h00;
RAM[16'h7744] = 8'h00;
RAM[16'h7745] = 8'h00;
RAM[16'h7746] = 8'h00;
RAM[16'h7747] = 8'h00;
RAM[16'h7748] = 8'h00;
RAM[16'h7749] = 8'h00;
RAM[16'h774A] = 8'h00;
RAM[16'h774B] = 8'h00;
RAM[16'h774C] = 8'h00;
RAM[16'h774D] = 8'h00;
RAM[16'h774E] = 8'h00;
RAM[16'h774F] = 8'h00;
RAM[16'h7750] = 8'h00;
RAM[16'h7751] = 8'h00;
RAM[16'h7752] = 8'h00;
RAM[16'h7753] = 8'h00;
RAM[16'h7754] = 8'h00;
RAM[16'h7755] = 8'h00;
RAM[16'h7756] = 8'h00;
RAM[16'h7757] = 8'h00;
RAM[16'h7758] = 8'h00;
RAM[16'h7759] = 8'h00;
RAM[16'h775A] = 8'h00;
RAM[16'h775B] = 8'h00;
RAM[16'h775C] = 8'h00;
RAM[16'h775D] = 8'h00;
RAM[16'h775E] = 8'h00;
RAM[16'h775F] = 8'h00;
RAM[16'h7760] = 8'h00;
RAM[16'h7761] = 8'h00;
RAM[16'h7762] = 8'h00;
RAM[16'h7763] = 8'h00;
RAM[16'h7764] = 8'h00;
RAM[16'h7765] = 8'h00;
RAM[16'h7766] = 8'h00;
RAM[16'h7767] = 8'h00;
RAM[16'h7768] = 8'h00;
RAM[16'h7769] = 8'h00;
RAM[16'h776A] = 8'h00;
RAM[16'h776B] = 8'h00;
RAM[16'h776C] = 8'h00;
RAM[16'h776D] = 8'h00;
RAM[16'h776E] = 8'h00;
RAM[16'h776F] = 8'h00;
RAM[16'h7770] = 8'h00;
RAM[16'h7771] = 8'h00;
RAM[16'h7772] = 8'h00;
RAM[16'h7773] = 8'h00;
RAM[16'h7774] = 8'h00;
RAM[16'h7775] = 8'h00;
RAM[16'h7776] = 8'h00;
RAM[16'h7777] = 8'h00;
RAM[16'h7778] = 8'h00;
RAM[16'h7779] = 8'h00;
RAM[16'h777A] = 8'h00;
RAM[16'h777B] = 8'h00;
RAM[16'h777C] = 8'h00;
RAM[16'h777D] = 8'h00;
RAM[16'h777E] = 8'h00;
RAM[16'h777F] = 8'h00;
RAM[16'h7780] = 8'h00;
RAM[16'h7781] = 8'h00;
RAM[16'h7782] = 8'h00;
RAM[16'h7783] = 8'h00;
RAM[16'h7784] = 8'h00;
RAM[16'h7785] = 8'h00;
RAM[16'h7786] = 8'h00;
RAM[16'h7787] = 8'h00;
RAM[16'h7788] = 8'h00;
RAM[16'h7789] = 8'h00;
RAM[16'h778A] = 8'h00;
RAM[16'h778B] = 8'h00;
RAM[16'h778C] = 8'h00;
RAM[16'h778D] = 8'h00;
RAM[16'h778E] = 8'h00;
RAM[16'h778F] = 8'h00;
RAM[16'h7790] = 8'h00;
RAM[16'h7791] = 8'h00;
RAM[16'h7792] = 8'h00;
RAM[16'h7793] = 8'h00;
RAM[16'h7794] = 8'h00;
RAM[16'h7795] = 8'h00;
RAM[16'h7796] = 8'h00;
RAM[16'h7797] = 8'h00;
RAM[16'h7798] = 8'h00;
RAM[16'h7799] = 8'h00;
RAM[16'h779A] = 8'h00;
RAM[16'h779B] = 8'h00;
RAM[16'h779C] = 8'h00;
RAM[16'h779D] = 8'h00;
RAM[16'h779E] = 8'h00;
RAM[16'h779F] = 8'h00;
RAM[16'h77A0] = 8'h00;
RAM[16'h77A1] = 8'h00;
RAM[16'h77A2] = 8'h00;
RAM[16'h77A3] = 8'h00;
RAM[16'h77A4] = 8'h00;
RAM[16'h77A5] = 8'h00;
RAM[16'h77A6] = 8'h00;
RAM[16'h77A7] = 8'h00;
RAM[16'h77A8] = 8'h00;
RAM[16'h77A9] = 8'h00;
RAM[16'h77AA] = 8'h00;
RAM[16'h77AB] = 8'h00;
RAM[16'h77AC] = 8'h00;
RAM[16'h77AD] = 8'h00;
RAM[16'h77AE] = 8'h00;
RAM[16'h77AF] = 8'h00;
RAM[16'h77B0] = 8'h00;
RAM[16'h77B1] = 8'h00;
RAM[16'h77B2] = 8'h00;
RAM[16'h77B3] = 8'h00;
RAM[16'h77B4] = 8'h00;
RAM[16'h77B5] = 8'h00;
RAM[16'h77B6] = 8'h00;
RAM[16'h77B7] = 8'h00;
RAM[16'h77B8] = 8'h00;
RAM[16'h77B9] = 8'h00;
RAM[16'h77BA] = 8'h00;
RAM[16'h77BB] = 8'h00;
RAM[16'h77BC] = 8'h00;
RAM[16'h77BD] = 8'h00;
RAM[16'h77BE] = 8'h00;
RAM[16'h77BF] = 8'h00;
RAM[16'h77C0] = 8'h00;
RAM[16'h77C1] = 8'h00;
RAM[16'h77C2] = 8'h00;
RAM[16'h77C3] = 8'h00;
RAM[16'h77C4] = 8'h00;
RAM[16'h77C5] = 8'h00;
RAM[16'h77C6] = 8'h00;
RAM[16'h77C7] = 8'h00;
RAM[16'h77C8] = 8'h00;
RAM[16'h77C9] = 8'h00;
RAM[16'h77CA] = 8'h00;
RAM[16'h77CB] = 8'h00;
RAM[16'h77CC] = 8'h00;
RAM[16'h77CD] = 8'h00;
RAM[16'h77CE] = 8'h00;
RAM[16'h77CF] = 8'h00;
RAM[16'h77D0] = 8'h00;
RAM[16'h77D1] = 8'h00;
RAM[16'h77D2] = 8'h00;
RAM[16'h77D3] = 8'h00;
RAM[16'h77D4] = 8'h00;
RAM[16'h77D5] = 8'h00;
RAM[16'h77D6] = 8'h00;
RAM[16'h77D7] = 8'h00;
RAM[16'h77D8] = 8'h00;
RAM[16'h77D9] = 8'h00;
RAM[16'h77DA] = 8'h00;
RAM[16'h77DB] = 8'h00;
RAM[16'h77DC] = 8'h00;
RAM[16'h77DD] = 8'h00;
RAM[16'h77DE] = 8'h00;
RAM[16'h77DF] = 8'h00;
RAM[16'h77E0] = 8'h00;
RAM[16'h77E1] = 8'h00;
RAM[16'h77E2] = 8'h00;
RAM[16'h77E3] = 8'h00;
RAM[16'h77E4] = 8'h00;
RAM[16'h77E5] = 8'h00;
RAM[16'h77E6] = 8'h00;
RAM[16'h77E7] = 8'h00;
RAM[16'h77E8] = 8'h00;
RAM[16'h77E9] = 8'h00;
RAM[16'h77EA] = 8'h00;
RAM[16'h77EB] = 8'h00;
RAM[16'h77EC] = 8'h00;
RAM[16'h77ED] = 8'h00;
RAM[16'h77EE] = 8'h00;
RAM[16'h77EF] = 8'h00;
RAM[16'h77F0] = 8'h00;
RAM[16'h77F1] = 8'h00;
RAM[16'h77F2] = 8'h00;
RAM[16'h77F3] = 8'h00;
RAM[16'h77F4] = 8'h00;
RAM[16'h77F5] = 8'h00;
RAM[16'h77F6] = 8'h00;
RAM[16'h77F7] = 8'h00;
RAM[16'h77F8] = 8'h00;
RAM[16'h77F9] = 8'h00;
RAM[16'h77FA] = 8'h00;
RAM[16'h77FB] = 8'h00;
RAM[16'h77FC] = 8'h00;
RAM[16'h77FD] = 8'h00;
RAM[16'h77FE] = 8'h00;
RAM[16'h77FF] = 8'h00;
RAM[16'h7800] = 8'h00;
RAM[16'h7801] = 8'h00;
RAM[16'h7802] = 8'h00;
RAM[16'h7803] = 8'h00;
RAM[16'h7804] = 8'h00;
RAM[16'h7805] = 8'h00;
RAM[16'h7806] = 8'h00;
RAM[16'h7807] = 8'h00;
RAM[16'h7808] = 8'h00;
RAM[16'h7809] = 8'h00;
RAM[16'h780A] = 8'h00;
RAM[16'h780B] = 8'h00;
RAM[16'h780C] = 8'h00;
RAM[16'h780D] = 8'h00;
RAM[16'h780E] = 8'h00;
RAM[16'h780F] = 8'h00;
RAM[16'h7810] = 8'h00;
RAM[16'h7811] = 8'h00;
RAM[16'h7812] = 8'h00;
RAM[16'h7813] = 8'h00;
RAM[16'h7814] = 8'h00;
RAM[16'h7815] = 8'h00;
RAM[16'h7816] = 8'h00;
RAM[16'h7817] = 8'h00;
RAM[16'h7818] = 8'h00;
RAM[16'h7819] = 8'h00;
RAM[16'h781A] = 8'h00;
RAM[16'h781B] = 8'h00;
RAM[16'h781C] = 8'h00;
RAM[16'h781D] = 8'h00;
RAM[16'h781E] = 8'h00;
RAM[16'h781F] = 8'h00;
RAM[16'h7820] = 8'h00;
RAM[16'h7821] = 8'h00;
RAM[16'h7822] = 8'h00;
RAM[16'h7823] = 8'h00;
RAM[16'h7824] = 8'h00;
RAM[16'h7825] = 8'h00;
RAM[16'h7826] = 8'h00;
RAM[16'h7827] = 8'h00;
RAM[16'h7828] = 8'h00;
RAM[16'h7829] = 8'h00;
RAM[16'h782A] = 8'h00;
RAM[16'h782B] = 8'h00;
RAM[16'h782C] = 8'h00;
RAM[16'h782D] = 8'h00;
RAM[16'h782E] = 8'h00;
RAM[16'h782F] = 8'h00;
RAM[16'h7830] = 8'h00;
RAM[16'h7831] = 8'h00;
RAM[16'h7832] = 8'h00;
RAM[16'h7833] = 8'h00;
RAM[16'h7834] = 8'h00;
RAM[16'h7835] = 8'h00;
RAM[16'h7836] = 8'h00;
RAM[16'h7837] = 8'h00;
RAM[16'h7838] = 8'h00;
RAM[16'h7839] = 8'h00;
RAM[16'h783A] = 8'h00;
RAM[16'h783B] = 8'h00;
RAM[16'h783C] = 8'h00;
RAM[16'h783D] = 8'h00;
RAM[16'h783E] = 8'h00;
RAM[16'h783F] = 8'h00;
RAM[16'h7840] = 8'h00;
RAM[16'h7841] = 8'h00;
RAM[16'h7842] = 8'h00;
RAM[16'h7843] = 8'h00;
RAM[16'h7844] = 8'h00;
RAM[16'h7845] = 8'h00;
RAM[16'h7846] = 8'h00;
RAM[16'h7847] = 8'h00;
RAM[16'h7848] = 8'h00;
RAM[16'h7849] = 8'h00;
RAM[16'h784A] = 8'h00;
RAM[16'h784B] = 8'h00;
RAM[16'h784C] = 8'h00;
RAM[16'h784D] = 8'h00;
RAM[16'h784E] = 8'h00;
RAM[16'h784F] = 8'h00;
RAM[16'h7850] = 8'h00;
RAM[16'h7851] = 8'h00;
RAM[16'h7852] = 8'h00;
RAM[16'h7853] = 8'h00;
RAM[16'h7854] = 8'h00;
RAM[16'h7855] = 8'h00;
RAM[16'h7856] = 8'h00;
RAM[16'h7857] = 8'h00;
RAM[16'h7858] = 8'h00;
RAM[16'h7859] = 8'h00;
RAM[16'h785A] = 8'h00;
RAM[16'h785B] = 8'h00;
RAM[16'h785C] = 8'h00;
RAM[16'h785D] = 8'h00;
RAM[16'h785E] = 8'h00;
RAM[16'h785F] = 8'h00;
RAM[16'h7860] = 8'h00;
RAM[16'h7861] = 8'h00;
RAM[16'h7862] = 8'h00;
RAM[16'h7863] = 8'h00;
RAM[16'h7864] = 8'h00;
RAM[16'h7865] = 8'h00;
RAM[16'h7866] = 8'h00;
RAM[16'h7867] = 8'h00;
RAM[16'h7868] = 8'h00;
RAM[16'h7869] = 8'h00;
RAM[16'h786A] = 8'h00;
RAM[16'h786B] = 8'h00;
RAM[16'h786C] = 8'h00;
RAM[16'h786D] = 8'h00;
RAM[16'h786E] = 8'h00;
RAM[16'h786F] = 8'h00;
RAM[16'h7870] = 8'h00;
RAM[16'h7871] = 8'h00;
RAM[16'h7872] = 8'h00;
RAM[16'h7873] = 8'h00;
RAM[16'h7874] = 8'h00;
RAM[16'h7875] = 8'h00;
RAM[16'h7876] = 8'h00;
RAM[16'h7877] = 8'h00;
RAM[16'h7878] = 8'h00;
RAM[16'h7879] = 8'h00;
RAM[16'h787A] = 8'h00;
RAM[16'h787B] = 8'h00;
RAM[16'h787C] = 8'h00;
RAM[16'h787D] = 8'h00;
RAM[16'h787E] = 8'h00;
RAM[16'h787F] = 8'h00;
RAM[16'h7880] = 8'h00;
RAM[16'h7881] = 8'h00;
RAM[16'h7882] = 8'h00;
RAM[16'h7883] = 8'h00;
RAM[16'h7884] = 8'h00;
RAM[16'h7885] = 8'h00;
RAM[16'h7886] = 8'h00;
RAM[16'h7887] = 8'h00;
RAM[16'h7888] = 8'h00;
RAM[16'h7889] = 8'h00;
RAM[16'h788A] = 8'h00;
RAM[16'h788B] = 8'h00;
RAM[16'h788C] = 8'h00;
RAM[16'h788D] = 8'h00;
RAM[16'h788E] = 8'h00;
RAM[16'h788F] = 8'h00;
RAM[16'h7890] = 8'h00;
RAM[16'h7891] = 8'h00;
RAM[16'h7892] = 8'h00;
RAM[16'h7893] = 8'h00;
RAM[16'h7894] = 8'h00;
RAM[16'h7895] = 8'h00;
RAM[16'h7896] = 8'h00;
RAM[16'h7897] = 8'h00;
RAM[16'h7898] = 8'h00;
RAM[16'h7899] = 8'h00;
RAM[16'h789A] = 8'h00;
RAM[16'h789B] = 8'h00;
RAM[16'h789C] = 8'h00;
RAM[16'h789D] = 8'h00;
RAM[16'h789E] = 8'h00;
RAM[16'h789F] = 8'h00;
RAM[16'h78A0] = 8'h00;
RAM[16'h78A1] = 8'h00;
RAM[16'h78A2] = 8'h00;
RAM[16'h78A3] = 8'h00;
RAM[16'h78A4] = 8'h00;
RAM[16'h78A5] = 8'h00;
RAM[16'h78A6] = 8'h00;
RAM[16'h78A7] = 8'h00;
RAM[16'h78A8] = 8'h00;
RAM[16'h78A9] = 8'h00;
RAM[16'h78AA] = 8'h00;
RAM[16'h78AB] = 8'h00;
RAM[16'h78AC] = 8'h00;
RAM[16'h78AD] = 8'h00;
RAM[16'h78AE] = 8'h00;
RAM[16'h78AF] = 8'h00;
RAM[16'h78B0] = 8'h00;
RAM[16'h78B1] = 8'h00;
RAM[16'h78B2] = 8'h00;
RAM[16'h78B3] = 8'h00;
RAM[16'h78B4] = 8'h00;
RAM[16'h78B5] = 8'h00;
RAM[16'h78B6] = 8'h00;
RAM[16'h78B7] = 8'h00;
RAM[16'h78B8] = 8'h00;
RAM[16'h78B9] = 8'h00;
RAM[16'h78BA] = 8'h00;
RAM[16'h78BB] = 8'h00;
RAM[16'h78BC] = 8'h00;
RAM[16'h78BD] = 8'h00;
RAM[16'h78BE] = 8'h00;
RAM[16'h78BF] = 8'h00;
RAM[16'h78C0] = 8'h00;
RAM[16'h78C1] = 8'h00;
RAM[16'h78C2] = 8'h00;
RAM[16'h78C3] = 8'h00;
RAM[16'h78C4] = 8'h00;
RAM[16'h78C5] = 8'h00;
RAM[16'h78C6] = 8'h00;
RAM[16'h78C7] = 8'h00;
RAM[16'h78C8] = 8'h00;
RAM[16'h78C9] = 8'h00;
RAM[16'h78CA] = 8'h00;
RAM[16'h78CB] = 8'h00;
RAM[16'h78CC] = 8'h00;
RAM[16'h78CD] = 8'h00;
RAM[16'h78CE] = 8'h00;
RAM[16'h78CF] = 8'h00;
RAM[16'h78D0] = 8'h00;
RAM[16'h78D1] = 8'h00;
RAM[16'h78D2] = 8'h00;
RAM[16'h78D3] = 8'h00;
RAM[16'h78D4] = 8'h00;
RAM[16'h78D5] = 8'h00;
RAM[16'h78D6] = 8'h00;
RAM[16'h78D7] = 8'h00;
RAM[16'h78D8] = 8'h00;
RAM[16'h78D9] = 8'h00;
RAM[16'h78DA] = 8'h00;
RAM[16'h78DB] = 8'h00;
RAM[16'h78DC] = 8'h00;
RAM[16'h78DD] = 8'h00;
RAM[16'h78DE] = 8'h00;
RAM[16'h78DF] = 8'h00;
RAM[16'h78E0] = 8'h00;
RAM[16'h78E1] = 8'h00;
RAM[16'h78E2] = 8'h00;
RAM[16'h78E3] = 8'h00;
RAM[16'h78E4] = 8'h00;
RAM[16'h78E5] = 8'h00;
RAM[16'h78E6] = 8'h00;
RAM[16'h78E7] = 8'h00;
RAM[16'h78E8] = 8'h00;
RAM[16'h78E9] = 8'h00;
RAM[16'h78EA] = 8'h00;
RAM[16'h78EB] = 8'h00;
RAM[16'h78EC] = 8'h00;
RAM[16'h78ED] = 8'h00;
RAM[16'h78EE] = 8'h00;
RAM[16'h78EF] = 8'h00;
RAM[16'h78F0] = 8'h00;
RAM[16'h78F1] = 8'h00;
RAM[16'h78F2] = 8'h00;
RAM[16'h78F3] = 8'h00;
RAM[16'h78F4] = 8'h00;
RAM[16'h78F5] = 8'h00;
RAM[16'h78F6] = 8'h00;
RAM[16'h78F7] = 8'h00;
RAM[16'h78F8] = 8'h00;
RAM[16'h78F9] = 8'h00;
RAM[16'h78FA] = 8'h00;
RAM[16'h78FB] = 8'h00;
RAM[16'h78FC] = 8'h00;
RAM[16'h78FD] = 8'h00;
RAM[16'h78FE] = 8'h00;
RAM[16'h78FF] = 8'h00;
RAM[16'h7900] = 8'h00;
RAM[16'h7901] = 8'h00;
RAM[16'h7902] = 8'h00;
RAM[16'h7903] = 8'h00;
RAM[16'h7904] = 8'h00;
RAM[16'h7905] = 8'h00;
RAM[16'h7906] = 8'h00;
RAM[16'h7907] = 8'h00;
RAM[16'h7908] = 8'h00;
RAM[16'h7909] = 8'h00;
RAM[16'h790A] = 8'h00;
RAM[16'h790B] = 8'h00;
RAM[16'h790C] = 8'h00;
RAM[16'h790D] = 8'h00;
RAM[16'h790E] = 8'h00;
RAM[16'h790F] = 8'h00;
RAM[16'h7910] = 8'h00;
RAM[16'h7911] = 8'h00;
RAM[16'h7912] = 8'h00;
RAM[16'h7913] = 8'h00;
RAM[16'h7914] = 8'h00;
RAM[16'h7915] = 8'h00;
RAM[16'h7916] = 8'h00;
RAM[16'h7917] = 8'h00;
RAM[16'h7918] = 8'h00;
RAM[16'h7919] = 8'h00;
RAM[16'h791A] = 8'h00;
RAM[16'h791B] = 8'h00;
RAM[16'h791C] = 8'h00;
RAM[16'h791D] = 8'h00;
RAM[16'h791E] = 8'h00;
RAM[16'h791F] = 8'h00;
RAM[16'h7920] = 8'h00;
RAM[16'h7921] = 8'h00;
RAM[16'h7922] = 8'h00;
RAM[16'h7923] = 8'h00;
RAM[16'h7924] = 8'h00;
RAM[16'h7925] = 8'h00;
RAM[16'h7926] = 8'h00;
RAM[16'h7927] = 8'h00;
RAM[16'h7928] = 8'h00;
RAM[16'h7929] = 8'h00;
RAM[16'h792A] = 8'h00;
RAM[16'h792B] = 8'h00;
RAM[16'h792C] = 8'h00;
RAM[16'h792D] = 8'h00;
RAM[16'h792E] = 8'h00;
RAM[16'h792F] = 8'h00;
RAM[16'h7930] = 8'h00;
RAM[16'h7931] = 8'h00;
RAM[16'h7932] = 8'h00;
RAM[16'h7933] = 8'h00;
RAM[16'h7934] = 8'h00;
RAM[16'h7935] = 8'h00;
RAM[16'h7936] = 8'h00;
RAM[16'h7937] = 8'h00;
RAM[16'h7938] = 8'h00;
RAM[16'h7939] = 8'h00;
RAM[16'h793A] = 8'h00;
RAM[16'h793B] = 8'h00;
RAM[16'h793C] = 8'h00;
RAM[16'h793D] = 8'h00;
RAM[16'h793E] = 8'h00;
RAM[16'h793F] = 8'h00;
RAM[16'h7940] = 8'h00;
RAM[16'h7941] = 8'h00;
RAM[16'h7942] = 8'h00;
RAM[16'h7943] = 8'h00;
RAM[16'h7944] = 8'h00;
RAM[16'h7945] = 8'h00;
RAM[16'h7946] = 8'h00;
RAM[16'h7947] = 8'h00;
RAM[16'h7948] = 8'h00;
RAM[16'h7949] = 8'h00;
RAM[16'h794A] = 8'h00;
RAM[16'h794B] = 8'h00;
RAM[16'h794C] = 8'h00;
RAM[16'h794D] = 8'h00;
RAM[16'h794E] = 8'h00;
RAM[16'h794F] = 8'h00;
RAM[16'h7950] = 8'h00;
RAM[16'h7951] = 8'h00;
RAM[16'h7952] = 8'h00;
RAM[16'h7953] = 8'h00;
RAM[16'h7954] = 8'h00;
RAM[16'h7955] = 8'h00;
RAM[16'h7956] = 8'h00;
RAM[16'h7957] = 8'h00;
RAM[16'h7958] = 8'h00;
RAM[16'h7959] = 8'h00;
RAM[16'h795A] = 8'h00;
RAM[16'h795B] = 8'h00;
RAM[16'h795C] = 8'h00;
RAM[16'h795D] = 8'h00;
RAM[16'h795E] = 8'h00;
RAM[16'h795F] = 8'h00;
RAM[16'h7960] = 8'h00;
RAM[16'h7961] = 8'h00;
RAM[16'h7962] = 8'h00;
RAM[16'h7963] = 8'h00;
RAM[16'h7964] = 8'h00;
RAM[16'h7965] = 8'h00;
RAM[16'h7966] = 8'h00;
RAM[16'h7967] = 8'h00;
RAM[16'h7968] = 8'h00;
RAM[16'h7969] = 8'h00;
RAM[16'h796A] = 8'h00;
RAM[16'h796B] = 8'h00;
RAM[16'h796C] = 8'h00;
RAM[16'h796D] = 8'h00;
RAM[16'h796E] = 8'h00;
RAM[16'h796F] = 8'h00;
RAM[16'h7970] = 8'h00;
RAM[16'h7971] = 8'h00;
RAM[16'h7972] = 8'h00;
RAM[16'h7973] = 8'h00;
RAM[16'h7974] = 8'h00;
RAM[16'h7975] = 8'h00;
RAM[16'h7976] = 8'h00;
RAM[16'h7977] = 8'h00;
RAM[16'h7978] = 8'h00;
RAM[16'h7979] = 8'h00;
RAM[16'h797A] = 8'h00;
RAM[16'h797B] = 8'h00;
RAM[16'h797C] = 8'h00;
RAM[16'h797D] = 8'h00;
RAM[16'h797E] = 8'h00;
RAM[16'h797F] = 8'h00;
RAM[16'h7980] = 8'h00;
RAM[16'h7981] = 8'h00;
RAM[16'h7982] = 8'h00;
RAM[16'h7983] = 8'h00;
RAM[16'h7984] = 8'h00;
RAM[16'h7985] = 8'h00;
RAM[16'h7986] = 8'h00;
RAM[16'h7987] = 8'h00;
RAM[16'h7988] = 8'h00;
RAM[16'h7989] = 8'h00;
RAM[16'h798A] = 8'h00;
RAM[16'h798B] = 8'h00;
RAM[16'h798C] = 8'h00;
RAM[16'h798D] = 8'h00;
RAM[16'h798E] = 8'h00;
RAM[16'h798F] = 8'h00;
RAM[16'h7990] = 8'h00;
RAM[16'h7991] = 8'h00;
RAM[16'h7992] = 8'h00;
RAM[16'h7993] = 8'h00;
RAM[16'h7994] = 8'h00;
RAM[16'h7995] = 8'h00;
RAM[16'h7996] = 8'h00;
RAM[16'h7997] = 8'h00;
RAM[16'h7998] = 8'h00;
RAM[16'h7999] = 8'h00;
RAM[16'h799A] = 8'h00;
RAM[16'h799B] = 8'h00;
RAM[16'h799C] = 8'h00;
RAM[16'h799D] = 8'h00;
RAM[16'h799E] = 8'h00;
RAM[16'h799F] = 8'h00;
RAM[16'h79A0] = 8'h00;
RAM[16'h79A1] = 8'h00;
RAM[16'h79A2] = 8'h00;
RAM[16'h79A3] = 8'h00;
RAM[16'h79A4] = 8'h00;
RAM[16'h79A5] = 8'h00;
RAM[16'h79A6] = 8'h00;
RAM[16'h79A7] = 8'h00;
RAM[16'h79A8] = 8'h00;
RAM[16'h79A9] = 8'h00;
RAM[16'h79AA] = 8'h00;
RAM[16'h79AB] = 8'h00;
RAM[16'h79AC] = 8'h00;
RAM[16'h79AD] = 8'h00;
RAM[16'h79AE] = 8'h00;
RAM[16'h79AF] = 8'h00;
RAM[16'h79B0] = 8'h00;
RAM[16'h79B1] = 8'h00;
RAM[16'h79B2] = 8'h00;
RAM[16'h79B3] = 8'h00;
RAM[16'h79B4] = 8'h00;
RAM[16'h79B5] = 8'h00;
RAM[16'h79B6] = 8'h00;
RAM[16'h79B7] = 8'h00;
RAM[16'h79B8] = 8'h00;
RAM[16'h79B9] = 8'h00;
RAM[16'h79BA] = 8'h00;
RAM[16'h79BB] = 8'h00;
RAM[16'h79BC] = 8'h00;
RAM[16'h79BD] = 8'h00;
RAM[16'h79BE] = 8'h00;
RAM[16'h79BF] = 8'h00;
RAM[16'h79C0] = 8'h00;
RAM[16'h79C1] = 8'h00;
RAM[16'h79C2] = 8'h00;
RAM[16'h79C3] = 8'h00;
RAM[16'h79C4] = 8'h00;
RAM[16'h79C5] = 8'h00;
RAM[16'h79C6] = 8'h00;
RAM[16'h79C7] = 8'h00;
RAM[16'h79C8] = 8'h00;
RAM[16'h79C9] = 8'h00;
RAM[16'h79CA] = 8'h00;
RAM[16'h79CB] = 8'h00;
RAM[16'h79CC] = 8'h00;
RAM[16'h79CD] = 8'h00;
RAM[16'h79CE] = 8'h00;
RAM[16'h79CF] = 8'h00;
RAM[16'h79D0] = 8'h00;
RAM[16'h79D1] = 8'h00;
RAM[16'h79D2] = 8'h00;
RAM[16'h79D3] = 8'h00;
RAM[16'h79D4] = 8'h00;
RAM[16'h79D5] = 8'h00;
RAM[16'h79D6] = 8'h00;
RAM[16'h79D7] = 8'h00;
RAM[16'h79D8] = 8'h00;
RAM[16'h79D9] = 8'h00;
RAM[16'h79DA] = 8'h00;
RAM[16'h79DB] = 8'h00;
RAM[16'h79DC] = 8'h00;
RAM[16'h79DD] = 8'h00;
RAM[16'h79DE] = 8'h00;
RAM[16'h79DF] = 8'h00;
RAM[16'h79E0] = 8'h00;
RAM[16'h79E1] = 8'h00;
RAM[16'h79E2] = 8'h00;
RAM[16'h79E3] = 8'h00;
RAM[16'h79E4] = 8'h00;
RAM[16'h79E5] = 8'h00;
RAM[16'h79E6] = 8'h00;
RAM[16'h79E7] = 8'h00;
RAM[16'h79E8] = 8'h00;
RAM[16'h79E9] = 8'h00;
RAM[16'h79EA] = 8'h00;
RAM[16'h79EB] = 8'h00;
RAM[16'h79EC] = 8'h00;
RAM[16'h79ED] = 8'h00;
RAM[16'h79EE] = 8'h00;
RAM[16'h79EF] = 8'h00;
RAM[16'h79F0] = 8'h00;
RAM[16'h79F1] = 8'h00;
RAM[16'h79F2] = 8'h00;
RAM[16'h79F3] = 8'h00;
RAM[16'h79F4] = 8'h00;
RAM[16'h79F5] = 8'h00;
RAM[16'h79F6] = 8'h00;
RAM[16'h79F7] = 8'h00;
RAM[16'h79F8] = 8'h00;
RAM[16'h79F9] = 8'h00;
RAM[16'h79FA] = 8'h00;
RAM[16'h79FB] = 8'h00;
RAM[16'h79FC] = 8'h00;
RAM[16'h79FD] = 8'h00;
RAM[16'h79FE] = 8'h00;
RAM[16'h79FF] = 8'h00;
RAM[16'h7A00] = 8'h00;
RAM[16'h7A01] = 8'h00;
RAM[16'h7A02] = 8'h00;
RAM[16'h7A03] = 8'h00;
RAM[16'h7A04] = 8'h00;
RAM[16'h7A05] = 8'h00;
RAM[16'h7A06] = 8'h00;
RAM[16'h7A07] = 8'h00;
RAM[16'h7A08] = 8'h00;
RAM[16'h7A09] = 8'h00;
RAM[16'h7A0A] = 8'h00;
RAM[16'h7A0B] = 8'h00;
RAM[16'h7A0C] = 8'h00;
RAM[16'h7A0D] = 8'h00;
RAM[16'h7A0E] = 8'h00;
RAM[16'h7A0F] = 8'h00;
RAM[16'h7A10] = 8'h00;
RAM[16'h7A11] = 8'h00;
RAM[16'h7A12] = 8'h00;
RAM[16'h7A13] = 8'h00;
RAM[16'h7A14] = 8'h00;
RAM[16'h7A15] = 8'h00;
RAM[16'h7A16] = 8'h00;
RAM[16'h7A17] = 8'h00;
RAM[16'h7A18] = 8'h00;
RAM[16'h7A19] = 8'h00;
RAM[16'h7A1A] = 8'h00;
RAM[16'h7A1B] = 8'h00;
RAM[16'h7A1C] = 8'h00;
RAM[16'h7A1D] = 8'h00;
RAM[16'h7A1E] = 8'h00;
RAM[16'h7A1F] = 8'h00;
RAM[16'h7A20] = 8'h00;
RAM[16'h7A21] = 8'h00;
RAM[16'h7A22] = 8'h00;
RAM[16'h7A23] = 8'h00;
RAM[16'h7A24] = 8'h00;
RAM[16'h7A25] = 8'h00;
RAM[16'h7A26] = 8'h00;
RAM[16'h7A27] = 8'h00;
RAM[16'h7A28] = 8'h00;
RAM[16'h7A29] = 8'h00;
RAM[16'h7A2A] = 8'h00;
RAM[16'h7A2B] = 8'h00;
RAM[16'h7A2C] = 8'h00;
RAM[16'h7A2D] = 8'h00;
RAM[16'h7A2E] = 8'h00;
RAM[16'h7A2F] = 8'h00;
RAM[16'h7A30] = 8'h00;
RAM[16'h7A31] = 8'h00;
RAM[16'h7A32] = 8'h00;
RAM[16'h7A33] = 8'h00;
RAM[16'h7A34] = 8'h00;
RAM[16'h7A35] = 8'h00;
RAM[16'h7A36] = 8'h00;
RAM[16'h7A37] = 8'h00;
RAM[16'h7A38] = 8'h00;
RAM[16'h7A39] = 8'h00;
RAM[16'h7A3A] = 8'h00;
RAM[16'h7A3B] = 8'h00;
RAM[16'h7A3C] = 8'h00;
RAM[16'h7A3D] = 8'h00;
RAM[16'h7A3E] = 8'h00;
RAM[16'h7A3F] = 8'h00;
RAM[16'h7A40] = 8'h00;
RAM[16'h7A41] = 8'h00;
RAM[16'h7A42] = 8'h00;
RAM[16'h7A43] = 8'h00;
RAM[16'h7A44] = 8'h00;
RAM[16'h7A45] = 8'h00;
RAM[16'h7A46] = 8'h00;
RAM[16'h7A47] = 8'h00;
RAM[16'h7A48] = 8'h00;
RAM[16'h7A49] = 8'h00;
RAM[16'h7A4A] = 8'h00;
RAM[16'h7A4B] = 8'h00;
RAM[16'h7A4C] = 8'h00;
RAM[16'h7A4D] = 8'h00;
RAM[16'h7A4E] = 8'h00;
RAM[16'h7A4F] = 8'h00;
RAM[16'h7A50] = 8'h00;
RAM[16'h7A51] = 8'h00;
RAM[16'h7A52] = 8'h00;
RAM[16'h7A53] = 8'h00;
RAM[16'h7A54] = 8'h00;
RAM[16'h7A55] = 8'h00;
RAM[16'h7A56] = 8'h00;
RAM[16'h7A57] = 8'h00;
RAM[16'h7A58] = 8'h00;
RAM[16'h7A59] = 8'h00;
RAM[16'h7A5A] = 8'h00;
RAM[16'h7A5B] = 8'h00;
RAM[16'h7A5C] = 8'h00;
RAM[16'h7A5D] = 8'h00;
RAM[16'h7A5E] = 8'h00;
RAM[16'h7A5F] = 8'h00;
RAM[16'h7A60] = 8'h00;
RAM[16'h7A61] = 8'h00;
RAM[16'h7A62] = 8'h00;
RAM[16'h7A63] = 8'h00;
RAM[16'h7A64] = 8'h00;
RAM[16'h7A65] = 8'h00;
RAM[16'h7A66] = 8'h00;
RAM[16'h7A67] = 8'h00;
RAM[16'h7A68] = 8'h00;
RAM[16'h7A69] = 8'h00;
RAM[16'h7A6A] = 8'h00;
RAM[16'h7A6B] = 8'h00;
RAM[16'h7A6C] = 8'h00;
RAM[16'h7A6D] = 8'h00;
RAM[16'h7A6E] = 8'h00;
RAM[16'h7A6F] = 8'h00;
RAM[16'h7A70] = 8'h00;
RAM[16'h7A71] = 8'h00;
RAM[16'h7A72] = 8'h00;
RAM[16'h7A73] = 8'h00;
RAM[16'h7A74] = 8'h00;
RAM[16'h7A75] = 8'h00;
RAM[16'h7A76] = 8'h00;
RAM[16'h7A77] = 8'h00;
RAM[16'h7A78] = 8'h00;
RAM[16'h7A79] = 8'h00;
RAM[16'h7A7A] = 8'h00;
RAM[16'h7A7B] = 8'h00;
RAM[16'h7A7C] = 8'h00;
RAM[16'h7A7D] = 8'h00;
RAM[16'h7A7E] = 8'h00;
RAM[16'h7A7F] = 8'h00;
RAM[16'h7A80] = 8'h00;
RAM[16'h7A81] = 8'h00;
RAM[16'h7A82] = 8'h00;
RAM[16'h7A83] = 8'h00;
RAM[16'h7A84] = 8'h00;
RAM[16'h7A85] = 8'h00;
RAM[16'h7A86] = 8'h00;
RAM[16'h7A87] = 8'h00;
RAM[16'h7A88] = 8'h00;
RAM[16'h7A89] = 8'h00;
RAM[16'h7A8A] = 8'h00;
RAM[16'h7A8B] = 8'h00;
RAM[16'h7A8C] = 8'h00;
RAM[16'h7A8D] = 8'h00;
RAM[16'h7A8E] = 8'h00;
RAM[16'h7A8F] = 8'h00;
RAM[16'h7A90] = 8'h00;
RAM[16'h7A91] = 8'h00;
RAM[16'h7A92] = 8'h00;
RAM[16'h7A93] = 8'h00;
RAM[16'h7A94] = 8'h00;
RAM[16'h7A95] = 8'h00;
RAM[16'h7A96] = 8'h00;
RAM[16'h7A97] = 8'h00;
RAM[16'h7A98] = 8'h00;
RAM[16'h7A99] = 8'h00;
RAM[16'h7A9A] = 8'h00;
RAM[16'h7A9B] = 8'h00;
RAM[16'h7A9C] = 8'h00;
RAM[16'h7A9D] = 8'h00;
RAM[16'h7A9E] = 8'h00;
RAM[16'h7A9F] = 8'h00;
RAM[16'h7AA0] = 8'h00;
RAM[16'h7AA1] = 8'h00;
RAM[16'h7AA2] = 8'h00;
RAM[16'h7AA3] = 8'h00;
RAM[16'h7AA4] = 8'h00;
RAM[16'h7AA5] = 8'h00;
RAM[16'h7AA6] = 8'h00;
RAM[16'h7AA7] = 8'h00;
RAM[16'h7AA8] = 8'h00;
RAM[16'h7AA9] = 8'h00;
RAM[16'h7AAA] = 8'h00;
RAM[16'h7AAB] = 8'h00;
RAM[16'h7AAC] = 8'h00;
RAM[16'h7AAD] = 8'h00;
RAM[16'h7AAE] = 8'h00;
RAM[16'h7AAF] = 8'h00;
RAM[16'h7AB0] = 8'h00;
RAM[16'h7AB1] = 8'h00;
RAM[16'h7AB2] = 8'h00;
RAM[16'h7AB3] = 8'h00;
RAM[16'h7AB4] = 8'h00;
RAM[16'h7AB5] = 8'h00;
RAM[16'h7AB6] = 8'h00;
RAM[16'h7AB7] = 8'h00;
RAM[16'h7AB8] = 8'h00;
RAM[16'h7AB9] = 8'h00;
RAM[16'h7ABA] = 8'h00;
RAM[16'h7ABB] = 8'h00;
RAM[16'h7ABC] = 8'h00;
RAM[16'h7ABD] = 8'h00;
RAM[16'h7ABE] = 8'h00;
RAM[16'h7ABF] = 8'h00;
RAM[16'h7AC0] = 8'h00;
RAM[16'h7AC1] = 8'h00;
RAM[16'h7AC2] = 8'h00;
RAM[16'h7AC3] = 8'h00;
RAM[16'h7AC4] = 8'h00;
RAM[16'h7AC5] = 8'h00;
RAM[16'h7AC6] = 8'h00;
RAM[16'h7AC7] = 8'h00;
RAM[16'h7AC8] = 8'h00;
RAM[16'h7AC9] = 8'h00;
RAM[16'h7ACA] = 8'h00;
RAM[16'h7ACB] = 8'h00;
RAM[16'h7ACC] = 8'h00;
RAM[16'h7ACD] = 8'h00;
RAM[16'h7ACE] = 8'h00;
RAM[16'h7ACF] = 8'h00;
RAM[16'h7AD0] = 8'h00;
RAM[16'h7AD1] = 8'h00;
RAM[16'h7AD2] = 8'h00;
RAM[16'h7AD3] = 8'h00;
RAM[16'h7AD4] = 8'h00;
RAM[16'h7AD5] = 8'h00;
RAM[16'h7AD6] = 8'h00;
RAM[16'h7AD7] = 8'h00;
RAM[16'h7AD8] = 8'h00;
RAM[16'h7AD9] = 8'h00;
RAM[16'h7ADA] = 8'h00;
RAM[16'h7ADB] = 8'h00;
RAM[16'h7ADC] = 8'h00;
RAM[16'h7ADD] = 8'h00;
RAM[16'h7ADE] = 8'h00;
RAM[16'h7ADF] = 8'h00;
RAM[16'h7AE0] = 8'h00;
RAM[16'h7AE1] = 8'h00;
RAM[16'h7AE2] = 8'h00;
RAM[16'h7AE3] = 8'h00;
RAM[16'h7AE4] = 8'h00;
RAM[16'h7AE5] = 8'h00;
RAM[16'h7AE6] = 8'h00;
RAM[16'h7AE7] = 8'h00;
RAM[16'h7AE8] = 8'h00;
RAM[16'h7AE9] = 8'h00;
RAM[16'h7AEA] = 8'h00;
RAM[16'h7AEB] = 8'h00;
RAM[16'h7AEC] = 8'h00;
RAM[16'h7AED] = 8'h00;
RAM[16'h7AEE] = 8'h00;
RAM[16'h7AEF] = 8'h00;
RAM[16'h7AF0] = 8'h00;
RAM[16'h7AF1] = 8'h00;
RAM[16'h7AF2] = 8'h00;
RAM[16'h7AF3] = 8'h00;
RAM[16'h7AF4] = 8'h00;
RAM[16'h7AF5] = 8'h00;
RAM[16'h7AF6] = 8'h00;
RAM[16'h7AF7] = 8'h00;
RAM[16'h7AF8] = 8'h00;
RAM[16'h7AF9] = 8'h00;
RAM[16'h7AFA] = 8'h00;
RAM[16'h7AFB] = 8'h00;
RAM[16'h7AFC] = 8'h00;
RAM[16'h7AFD] = 8'h00;
RAM[16'h7AFE] = 8'h00;
RAM[16'h7AFF] = 8'h00;
RAM[16'h7B00] = 8'h00;
RAM[16'h7B01] = 8'h00;
RAM[16'h7B02] = 8'h00;
RAM[16'h7B03] = 8'h00;
RAM[16'h7B04] = 8'h00;
RAM[16'h7B05] = 8'h00;
RAM[16'h7B06] = 8'h00;
RAM[16'h7B07] = 8'h00;
RAM[16'h7B08] = 8'h00;
RAM[16'h7B09] = 8'h00;
RAM[16'h7B0A] = 8'h00;
RAM[16'h7B0B] = 8'h00;
RAM[16'h7B0C] = 8'h00;
RAM[16'h7B0D] = 8'h00;
RAM[16'h7B0E] = 8'h00;
RAM[16'h7B0F] = 8'h00;
RAM[16'h7B10] = 8'h00;
RAM[16'h7B11] = 8'h00;
RAM[16'h7B12] = 8'h00;
RAM[16'h7B13] = 8'h00;
RAM[16'h7B14] = 8'h00;
RAM[16'h7B15] = 8'h00;
RAM[16'h7B16] = 8'h00;
RAM[16'h7B17] = 8'h00;
RAM[16'h7B18] = 8'h00;
RAM[16'h7B19] = 8'h00;
RAM[16'h7B1A] = 8'h00;
RAM[16'h7B1B] = 8'h00;
RAM[16'h7B1C] = 8'h00;
RAM[16'h7B1D] = 8'h00;
RAM[16'h7B1E] = 8'h00;
RAM[16'h7B1F] = 8'h00;
RAM[16'h7B20] = 8'h00;
RAM[16'h7B21] = 8'h00;
RAM[16'h7B22] = 8'h00;
RAM[16'h7B23] = 8'h00;
RAM[16'h7B24] = 8'h00;
RAM[16'h7B25] = 8'h00;
RAM[16'h7B26] = 8'h00;
RAM[16'h7B27] = 8'h00;
RAM[16'h7B28] = 8'h00;
RAM[16'h7B29] = 8'h00;
RAM[16'h7B2A] = 8'h00;
RAM[16'h7B2B] = 8'h00;
RAM[16'h7B2C] = 8'h00;
RAM[16'h7B2D] = 8'h00;
RAM[16'h7B2E] = 8'h00;
RAM[16'h7B2F] = 8'h00;
RAM[16'h7B30] = 8'h00;
RAM[16'h7B31] = 8'h00;
RAM[16'h7B32] = 8'h00;
RAM[16'h7B33] = 8'h00;
RAM[16'h7B34] = 8'h00;
RAM[16'h7B35] = 8'h00;
RAM[16'h7B36] = 8'h00;
RAM[16'h7B37] = 8'h00;
RAM[16'h7B38] = 8'h00;
RAM[16'h7B39] = 8'h00;
RAM[16'h7B3A] = 8'h00;
RAM[16'h7B3B] = 8'h00;
RAM[16'h7B3C] = 8'h00;
RAM[16'h7B3D] = 8'h00;
RAM[16'h7B3E] = 8'h00;
RAM[16'h7B3F] = 8'h00;
RAM[16'h7B40] = 8'h00;
RAM[16'h7B41] = 8'h00;
RAM[16'h7B42] = 8'h00;
RAM[16'h7B43] = 8'h00;
RAM[16'h7B44] = 8'h00;
RAM[16'h7B45] = 8'h00;
RAM[16'h7B46] = 8'h00;
RAM[16'h7B47] = 8'h00;
RAM[16'h7B48] = 8'h00;
RAM[16'h7B49] = 8'h00;
RAM[16'h7B4A] = 8'h00;
RAM[16'h7B4B] = 8'h00;
RAM[16'h7B4C] = 8'h00;
RAM[16'h7B4D] = 8'h00;
RAM[16'h7B4E] = 8'h00;
RAM[16'h7B4F] = 8'h00;
RAM[16'h7B50] = 8'h00;
RAM[16'h7B51] = 8'h00;
RAM[16'h7B52] = 8'h00;
RAM[16'h7B53] = 8'h00;
RAM[16'h7B54] = 8'h00;
RAM[16'h7B55] = 8'h00;
RAM[16'h7B56] = 8'h00;
RAM[16'h7B57] = 8'h00;
RAM[16'h7B58] = 8'h00;
RAM[16'h7B59] = 8'h00;
RAM[16'h7B5A] = 8'h00;
RAM[16'h7B5B] = 8'h00;
RAM[16'h7B5C] = 8'h00;
RAM[16'h7B5D] = 8'h00;
RAM[16'h7B5E] = 8'h00;
RAM[16'h7B5F] = 8'h00;
RAM[16'h7B60] = 8'h00;
RAM[16'h7B61] = 8'h00;
RAM[16'h7B62] = 8'h00;
RAM[16'h7B63] = 8'h00;
RAM[16'h7B64] = 8'h00;
RAM[16'h7B65] = 8'h00;
RAM[16'h7B66] = 8'h00;
RAM[16'h7B67] = 8'h00;
RAM[16'h7B68] = 8'h00;
RAM[16'h7B69] = 8'h00;
RAM[16'h7B6A] = 8'h00;
RAM[16'h7B6B] = 8'h00;
RAM[16'h7B6C] = 8'h00;
RAM[16'h7B6D] = 8'h00;
RAM[16'h7B6E] = 8'h00;
RAM[16'h7B6F] = 8'h00;
RAM[16'h7B70] = 8'h00;
RAM[16'h7B71] = 8'h00;
RAM[16'h7B72] = 8'h00;
RAM[16'h7B73] = 8'h00;
RAM[16'h7B74] = 8'h00;
RAM[16'h7B75] = 8'h00;
RAM[16'h7B76] = 8'h00;
RAM[16'h7B77] = 8'h00;
RAM[16'h7B78] = 8'h00;
RAM[16'h7B79] = 8'h00;
RAM[16'h7B7A] = 8'h00;
RAM[16'h7B7B] = 8'h00;
RAM[16'h7B7C] = 8'h00;
RAM[16'h7B7D] = 8'h00;
RAM[16'h7B7E] = 8'h00;
RAM[16'h7B7F] = 8'h00;
RAM[16'h7B80] = 8'h00;
RAM[16'h7B81] = 8'h00;
RAM[16'h7B82] = 8'h00;
RAM[16'h7B83] = 8'h00;
RAM[16'h7B84] = 8'h00;
RAM[16'h7B85] = 8'h00;
RAM[16'h7B86] = 8'h00;
RAM[16'h7B87] = 8'h00;
RAM[16'h7B88] = 8'h00;
RAM[16'h7B89] = 8'h00;
RAM[16'h7B8A] = 8'h00;
RAM[16'h7B8B] = 8'h00;
RAM[16'h7B8C] = 8'h00;
RAM[16'h7B8D] = 8'h00;
RAM[16'h7B8E] = 8'h00;
RAM[16'h7B8F] = 8'h00;
RAM[16'h7B90] = 8'h00;
RAM[16'h7B91] = 8'h00;
RAM[16'h7B92] = 8'h00;
RAM[16'h7B93] = 8'h00;
RAM[16'h7B94] = 8'h00;
RAM[16'h7B95] = 8'h00;
RAM[16'h7B96] = 8'h00;
RAM[16'h7B97] = 8'h00;
RAM[16'h7B98] = 8'h00;
RAM[16'h7B99] = 8'h00;
RAM[16'h7B9A] = 8'h00;
RAM[16'h7B9B] = 8'h00;
RAM[16'h7B9C] = 8'h00;
RAM[16'h7B9D] = 8'h00;
RAM[16'h7B9E] = 8'h00;
RAM[16'h7B9F] = 8'h00;
RAM[16'h7BA0] = 8'h00;
RAM[16'h7BA1] = 8'h00;
RAM[16'h7BA2] = 8'h00;
RAM[16'h7BA3] = 8'h00;
RAM[16'h7BA4] = 8'h00;
RAM[16'h7BA5] = 8'h00;
RAM[16'h7BA6] = 8'h00;
RAM[16'h7BA7] = 8'h00;
RAM[16'h7BA8] = 8'h00;
RAM[16'h7BA9] = 8'h00;
RAM[16'h7BAA] = 8'h00;
RAM[16'h7BAB] = 8'h00;
RAM[16'h7BAC] = 8'h00;
RAM[16'h7BAD] = 8'h00;
RAM[16'h7BAE] = 8'h00;
RAM[16'h7BAF] = 8'h00;
RAM[16'h7BB0] = 8'h00;
RAM[16'h7BB1] = 8'h00;
RAM[16'h7BB2] = 8'h00;
RAM[16'h7BB3] = 8'h00;
RAM[16'h7BB4] = 8'h00;
RAM[16'h7BB5] = 8'h00;
RAM[16'h7BB6] = 8'h00;
RAM[16'h7BB7] = 8'h00;
RAM[16'h7BB8] = 8'h00;
RAM[16'h7BB9] = 8'h00;
RAM[16'h7BBA] = 8'h00;
RAM[16'h7BBB] = 8'h00;
RAM[16'h7BBC] = 8'h00;
RAM[16'h7BBD] = 8'h00;
RAM[16'h7BBE] = 8'h00;
RAM[16'h7BBF] = 8'h00;
RAM[16'h7BC0] = 8'h00;
RAM[16'h7BC1] = 8'h00;
RAM[16'h7BC2] = 8'h00;
RAM[16'h7BC3] = 8'h00;
RAM[16'h7BC4] = 8'h00;
RAM[16'h7BC5] = 8'h00;
RAM[16'h7BC6] = 8'h00;
RAM[16'h7BC7] = 8'h00;
RAM[16'h7BC8] = 8'h00;
RAM[16'h7BC9] = 8'h00;
RAM[16'h7BCA] = 8'h00;
RAM[16'h7BCB] = 8'h00;
RAM[16'h7BCC] = 8'h00;
RAM[16'h7BCD] = 8'h00;
RAM[16'h7BCE] = 8'h00;
RAM[16'h7BCF] = 8'h00;
RAM[16'h7BD0] = 8'h00;
RAM[16'h7BD1] = 8'h00;
RAM[16'h7BD2] = 8'h00;
RAM[16'h7BD3] = 8'h00;
RAM[16'h7BD4] = 8'h00;
RAM[16'h7BD5] = 8'h00;
RAM[16'h7BD6] = 8'h00;
RAM[16'h7BD7] = 8'h00;
RAM[16'h7BD8] = 8'h00;
RAM[16'h7BD9] = 8'h00;
RAM[16'h7BDA] = 8'h00;
RAM[16'h7BDB] = 8'h00;
RAM[16'h7BDC] = 8'h00;
RAM[16'h7BDD] = 8'h00;
RAM[16'h7BDE] = 8'h00;
RAM[16'h7BDF] = 8'h00;
RAM[16'h7BE0] = 8'h00;
RAM[16'h7BE1] = 8'h00;
RAM[16'h7BE2] = 8'h00;
RAM[16'h7BE3] = 8'h00;
RAM[16'h7BE4] = 8'h00;
RAM[16'h7BE5] = 8'h00;
RAM[16'h7BE6] = 8'h00;
RAM[16'h7BE7] = 8'h00;
RAM[16'h7BE8] = 8'h00;
RAM[16'h7BE9] = 8'h00;
RAM[16'h7BEA] = 8'h00;
RAM[16'h7BEB] = 8'h00;
RAM[16'h7BEC] = 8'h00;
RAM[16'h7BED] = 8'h00;
RAM[16'h7BEE] = 8'h00;
RAM[16'h7BEF] = 8'h00;
RAM[16'h7BF0] = 8'h00;
RAM[16'h7BF1] = 8'h00;
RAM[16'h7BF2] = 8'h00;
RAM[16'h7BF3] = 8'h00;
RAM[16'h7BF4] = 8'h00;
RAM[16'h7BF5] = 8'h00;
RAM[16'h7BF6] = 8'h00;
RAM[16'h7BF7] = 8'h00;
RAM[16'h7BF8] = 8'h00;
RAM[16'h7BF9] = 8'h00;
RAM[16'h7BFA] = 8'h00;
RAM[16'h7BFB] = 8'h00;
RAM[16'h7BFC] = 8'h00;
RAM[16'h7BFD] = 8'h00;
RAM[16'h7BFE] = 8'h00;
RAM[16'h7BFF] = 8'h00;
RAM[16'h7C00] = 8'h00;
RAM[16'h7C01] = 8'h00;
RAM[16'h7C02] = 8'h00;
RAM[16'h7C03] = 8'h00;
RAM[16'h7C04] = 8'h00;
RAM[16'h7C05] = 8'h00;
RAM[16'h7C06] = 8'h00;
RAM[16'h7C07] = 8'h00;
RAM[16'h7C08] = 8'h00;
RAM[16'h7C09] = 8'h00;
RAM[16'h7C0A] = 8'h00;
RAM[16'h7C0B] = 8'h00;
RAM[16'h7C0C] = 8'h00;
RAM[16'h7C0D] = 8'h00;
RAM[16'h7C0E] = 8'h00;
RAM[16'h7C0F] = 8'h00;
RAM[16'h7C10] = 8'h00;
RAM[16'h7C11] = 8'h00;
RAM[16'h7C12] = 8'h00;
RAM[16'h7C13] = 8'h00;
RAM[16'h7C14] = 8'h00;
RAM[16'h7C15] = 8'h00;
RAM[16'h7C16] = 8'h00;
RAM[16'h7C17] = 8'h00;
RAM[16'h7C18] = 8'h00;
RAM[16'h7C19] = 8'h00;
RAM[16'h7C1A] = 8'h00;
RAM[16'h7C1B] = 8'h00;
RAM[16'h7C1C] = 8'h00;
RAM[16'h7C1D] = 8'h00;
RAM[16'h7C1E] = 8'h00;
RAM[16'h7C1F] = 8'h00;
RAM[16'h7C20] = 8'h00;
RAM[16'h7C21] = 8'h00;
RAM[16'h7C22] = 8'h00;
RAM[16'h7C23] = 8'h00;
RAM[16'h7C24] = 8'h00;
RAM[16'h7C25] = 8'h00;
RAM[16'h7C26] = 8'h00;
RAM[16'h7C27] = 8'h00;
RAM[16'h7C28] = 8'h00;
RAM[16'h7C29] = 8'h00;
RAM[16'h7C2A] = 8'h00;
RAM[16'h7C2B] = 8'h00;
RAM[16'h7C2C] = 8'h00;
RAM[16'h7C2D] = 8'h00;
RAM[16'h7C2E] = 8'h00;
RAM[16'h7C2F] = 8'h00;
RAM[16'h7C30] = 8'h00;
RAM[16'h7C31] = 8'h00;
RAM[16'h7C32] = 8'h00;
RAM[16'h7C33] = 8'h00;
RAM[16'h7C34] = 8'h00;
RAM[16'h7C35] = 8'h00;
RAM[16'h7C36] = 8'h00;
RAM[16'h7C37] = 8'h00;
RAM[16'h7C38] = 8'h00;
RAM[16'h7C39] = 8'h00;
RAM[16'h7C3A] = 8'h00;
RAM[16'h7C3B] = 8'h00;
RAM[16'h7C3C] = 8'h00;
RAM[16'h7C3D] = 8'h00;
RAM[16'h7C3E] = 8'h00;
RAM[16'h7C3F] = 8'h00;
RAM[16'h7C40] = 8'h00;
RAM[16'h7C41] = 8'h00;
RAM[16'h7C42] = 8'h00;
RAM[16'h7C43] = 8'h00;
RAM[16'h7C44] = 8'h00;
RAM[16'h7C45] = 8'h00;
RAM[16'h7C46] = 8'h00;
RAM[16'h7C47] = 8'h00;
RAM[16'h7C48] = 8'h00;
RAM[16'h7C49] = 8'h00;
RAM[16'h7C4A] = 8'h00;
RAM[16'h7C4B] = 8'h00;
RAM[16'h7C4C] = 8'h00;
RAM[16'h7C4D] = 8'h00;
RAM[16'h7C4E] = 8'h00;
RAM[16'h7C4F] = 8'h00;
RAM[16'h7C50] = 8'h00;
RAM[16'h7C51] = 8'h00;
RAM[16'h7C52] = 8'h00;
RAM[16'h7C53] = 8'h00;
RAM[16'h7C54] = 8'h00;
RAM[16'h7C55] = 8'h00;
RAM[16'h7C56] = 8'h00;
RAM[16'h7C57] = 8'h00;
RAM[16'h7C58] = 8'h00;
RAM[16'h7C59] = 8'h00;
RAM[16'h7C5A] = 8'h00;
RAM[16'h7C5B] = 8'h00;
RAM[16'h7C5C] = 8'h00;
RAM[16'h7C5D] = 8'h00;
RAM[16'h7C5E] = 8'h00;
RAM[16'h7C5F] = 8'h00;
RAM[16'h7C60] = 8'h00;
RAM[16'h7C61] = 8'h00;
RAM[16'h7C62] = 8'h00;
RAM[16'h7C63] = 8'h00;
RAM[16'h7C64] = 8'h00;
RAM[16'h7C65] = 8'h00;
RAM[16'h7C66] = 8'h00;
RAM[16'h7C67] = 8'h00;
RAM[16'h7C68] = 8'h00;
RAM[16'h7C69] = 8'h00;
RAM[16'h7C6A] = 8'h00;
RAM[16'h7C6B] = 8'h00;
RAM[16'h7C6C] = 8'h00;
RAM[16'h7C6D] = 8'h00;
RAM[16'h7C6E] = 8'h00;
RAM[16'h7C6F] = 8'h00;
RAM[16'h7C70] = 8'h00;
RAM[16'h7C71] = 8'h00;
RAM[16'h7C72] = 8'h00;
RAM[16'h7C73] = 8'h00;
RAM[16'h7C74] = 8'h00;
RAM[16'h7C75] = 8'h00;
RAM[16'h7C76] = 8'h00;
RAM[16'h7C77] = 8'h00;
RAM[16'h7C78] = 8'h00;
RAM[16'h7C79] = 8'h00;
RAM[16'h7C7A] = 8'h00;
RAM[16'h7C7B] = 8'h00;
RAM[16'h7C7C] = 8'h00;
RAM[16'h7C7D] = 8'h00;
RAM[16'h7C7E] = 8'h00;
RAM[16'h7C7F] = 8'h00;
RAM[16'h7C80] = 8'h00;
RAM[16'h7C81] = 8'h00;
RAM[16'h7C82] = 8'h00;
RAM[16'h7C83] = 8'h00;
RAM[16'h7C84] = 8'h00;
RAM[16'h7C85] = 8'h00;
RAM[16'h7C86] = 8'h00;
RAM[16'h7C87] = 8'h00;
RAM[16'h7C88] = 8'h00;
RAM[16'h7C89] = 8'h00;
RAM[16'h7C8A] = 8'h00;
RAM[16'h7C8B] = 8'h00;
RAM[16'h7C8C] = 8'h00;
RAM[16'h7C8D] = 8'h00;
RAM[16'h7C8E] = 8'h00;
RAM[16'h7C8F] = 8'h00;
RAM[16'h7C90] = 8'h00;
RAM[16'h7C91] = 8'h00;
RAM[16'h7C92] = 8'h00;
RAM[16'h7C93] = 8'h00;
RAM[16'h7C94] = 8'h00;
RAM[16'h7C95] = 8'h00;
RAM[16'h7C96] = 8'h00;
RAM[16'h7C97] = 8'h00;
RAM[16'h7C98] = 8'h00;
RAM[16'h7C99] = 8'h00;
RAM[16'h7C9A] = 8'h00;
RAM[16'h7C9B] = 8'h00;
RAM[16'h7C9C] = 8'h00;
RAM[16'h7C9D] = 8'h00;
RAM[16'h7C9E] = 8'h00;
RAM[16'h7C9F] = 8'h00;
RAM[16'h7CA0] = 8'h00;
RAM[16'h7CA1] = 8'h00;
RAM[16'h7CA2] = 8'h00;
RAM[16'h7CA3] = 8'h00;
RAM[16'h7CA4] = 8'h00;
RAM[16'h7CA5] = 8'h00;
RAM[16'h7CA6] = 8'h00;
RAM[16'h7CA7] = 8'h00;
RAM[16'h7CA8] = 8'h00;
RAM[16'h7CA9] = 8'h00;
RAM[16'h7CAA] = 8'h00;
RAM[16'h7CAB] = 8'h00;
RAM[16'h7CAC] = 8'h00;
RAM[16'h7CAD] = 8'h00;
RAM[16'h7CAE] = 8'h00;
RAM[16'h7CAF] = 8'h00;
RAM[16'h7CB0] = 8'h00;
RAM[16'h7CB1] = 8'h00;
RAM[16'h7CB2] = 8'h00;
RAM[16'h7CB3] = 8'h00;
RAM[16'h7CB4] = 8'h00;
RAM[16'h7CB5] = 8'h00;
RAM[16'h7CB6] = 8'h00;
RAM[16'h7CB7] = 8'h00;
RAM[16'h7CB8] = 8'h00;
RAM[16'h7CB9] = 8'h00;
RAM[16'h7CBA] = 8'h00;
RAM[16'h7CBB] = 8'h00;
RAM[16'h7CBC] = 8'h00;
RAM[16'h7CBD] = 8'h00;
RAM[16'h7CBE] = 8'h00;
RAM[16'h7CBF] = 8'h00;
RAM[16'h7CC0] = 8'h00;
RAM[16'h7CC1] = 8'h00;
RAM[16'h7CC2] = 8'h00;
RAM[16'h7CC3] = 8'h00;
RAM[16'h7CC4] = 8'h00;
RAM[16'h7CC5] = 8'h00;
RAM[16'h7CC6] = 8'h00;
RAM[16'h7CC7] = 8'h00;
RAM[16'h7CC8] = 8'h00;
RAM[16'h7CC9] = 8'h00;
RAM[16'h7CCA] = 8'h00;
RAM[16'h7CCB] = 8'h00;
RAM[16'h7CCC] = 8'h00;
RAM[16'h7CCD] = 8'h00;
RAM[16'h7CCE] = 8'h00;
RAM[16'h7CCF] = 8'h00;
RAM[16'h7CD0] = 8'h00;
RAM[16'h7CD1] = 8'h00;
RAM[16'h7CD2] = 8'h00;
RAM[16'h7CD3] = 8'h00;
RAM[16'h7CD4] = 8'h00;
RAM[16'h7CD5] = 8'h00;
RAM[16'h7CD6] = 8'h00;
RAM[16'h7CD7] = 8'h00;
RAM[16'h7CD8] = 8'h00;
RAM[16'h7CD9] = 8'h00;
RAM[16'h7CDA] = 8'h00;
RAM[16'h7CDB] = 8'h00;
RAM[16'h7CDC] = 8'h00;
RAM[16'h7CDD] = 8'h00;
RAM[16'h7CDE] = 8'h00;
RAM[16'h7CDF] = 8'h00;
RAM[16'h7CE0] = 8'h00;
RAM[16'h7CE1] = 8'h00;
RAM[16'h7CE2] = 8'h00;
RAM[16'h7CE3] = 8'h00;
RAM[16'h7CE4] = 8'h00;
RAM[16'h7CE5] = 8'h00;
RAM[16'h7CE6] = 8'h00;
RAM[16'h7CE7] = 8'h00;
RAM[16'h7CE8] = 8'h00;
RAM[16'h7CE9] = 8'h00;
RAM[16'h7CEA] = 8'h00;
RAM[16'h7CEB] = 8'h00;
RAM[16'h7CEC] = 8'h00;
RAM[16'h7CED] = 8'h00;
RAM[16'h7CEE] = 8'h00;
RAM[16'h7CEF] = 8'h00;
RAM[16'h7CF0] = 8'h00;
RAM[16'h7CF1] = 8'h00;
RAM[16'h7CF2] = 8'h00;
RAM[16'h7CF3] = 8'h00;
RAM[16'h7CF4] = 8'h00;
RAM[16'h7CF5] = 8'h00;
RAM[16'h7CF6] = 8'h00;
RAM[16'h7CF7] = 8'h00;
RAM[16'h7CF8] = 8'h00;
RAM[16'h7CF9] = 8'h00;
RAM[16'h7CFA] = 8'h00;
RAM[16'h7CFB] = 8'h00;
RAM[16'h7CFC] = 8'h00;
RAM[16'h7CFD] = 8'h00;
RAM[16'h7CFE] = 8'h00;
RAM[16'h7CFF] = 8'h00;
RAM[16'h7D00] = 8'h00;
RAM[16'h7D01] = 8'h00;
RAM[16'h7D02] = 8'h00;
RAM[16'h7D03] = 8'h00;
RAM[16'h7D04] = 8'h00;
RAM[16'h7D05] = 8'h00;
RAM[16'h7D06] = 8'h00;
RAM[16'h7D07] = 8'h00;
RAM[16'h7D08] = 8'h00;
RAM[16'h7D09] = 8'h00;
RAM[16'h7D0A] = 8'h00;
RAM[16'h7D0B] = 8'h00;
RAM[16'h7D0C] = 8'h00;
RAM[16'h7D0D] = 8'h00;
RAM[16'h7D0E] = 8'h00;
RAM[16'h7D0F] = 8'h00;
RAM[16'h7D10] = 8'h00;
RAM[16'h7D11] = 8'h00;
RAM[16'h7D12] = 8'h00;
RAM[16'h7D13] = 8'h00;
RAM[16'h7D14] = 8'h00;
RAM[16'h7D15] = 8'h00;
RAM[16'h7D16] = 8'h00;
RAM[16'h7D17] = 8'h00;
RAM[16'h7D18] = 8'h00;
RAM[16'h7D19] = 8'h00;
RAM[16'h7D1A] = 8'h00;
RAM[16'h7D1B] = 8'h00;
RAM[16'h7D1C] = 8'h00;
RAM[16'h7D1D] = 8'h00;
RAM[16'h7D1E] = 8'h00;
RAM[16'h7D1F] = 8'h00;
RAM[16'h7D20] = 8'h00;
RAM[16'h7D21] = 8'h00;
RAM[16'h7D22] = 8'h00;
RAM[16'h7D23] = 8'h00;
RAM[16'h7D24] = 8'h00;
RAM[16'h7D25] = 8'h00;
RAM[16'h7D26] = 8'h00;
RAM[16'h7D27] = 8'h00;
RAM[16'h7D28] = 8'h00;
RAM[16'h7D29] = 8'h00;
RAM[16'h7D2A] = 8'h00;
RAM[16'h7D2B] = 8'h00;
RAM[16'h7D2C] = 8'h00;
RAM[16'h7D2D] = 8'h00;
RAM[16'h7D2E] = 8'h00;
RAM[16'h7D2F] = 8'h00;
RAM[16'h7D30] = 8'h00;
RAM[16'h7D31] = 8'h00;
RAM[16'h7D32] = 8'h00;
RAM[16'h7D33] = 8'h00;
RAM[16'h7D34] = 8'h00;
RAM[16'h7D35] = 8'h00;
RAM[16'h7D36] = 8'h00;
RAM[16'h7D37] = 8'h00;
RAM[16'h7D38] = 8'h00;
RAM[16'h7D39] = 8'h00;
RAM[16'h7D3A] = 8'h00;
RAM[16'h7D3B] = 8'h00;
RAM[16'h7D3C] = 8'h00;
RAM[16'h7D3D] = 8'h00;
RAM[16'h7D3E] = 8'h00;
RAM[16'h7D3F] = 8'h00;
RAM[16'h7D40] = 8'h00;
RAM[16'h7D41] = 8'h00;
RAM[16'h7D42] = 8'h00;
RAM[16'h7D43] = 8'h00;
RAM[16'h7D44] = 8'h00;
RAM[16'h7D45] = 8'h00;
RAM[16'h7D46] = 8'h00;
RAM[16'h7D47] = 8'h00;
RAM[16'h7D48] = 8'h00;
RAM[16'h7D49] = 8'h00;
RAM[16'h7D4A] = 8'h00;
RAM[16'h7D4B] = 8'h00;
RAM[16'h7D4C] = 8'h00;
RAM[16'h7D4D] = 8'h00;
RAM[16'h7D4E] = 8'h00;
RAM[16'h7D4F] = 8'h00;
RAM[16'h7D50] = 8'h00;
RAM[16'h7D51] = 8'h00;
RAM[16'h7D52] = 8'h00;
RAM[16'h7D53] = 8'h00;
RAM[16'h7D54] = 8'h00;
RAM[16'h7D55] = 8'h00;
RAM[16'h7D56] = 8'h00;
RAM[16'h7D57] = 8'h00;
RAM[16'h7D58] = 8'h00;
RAM[16'h7D59] = 8'h00;
RAM[16'h7D5A] = 8'h00;
RAM[16'h7D5B] = 8'h00;
RAM[16'h7D5C] = 8'h00;
RAM[16'h7D5D] = 8'h00;
RAM[16'h7D5E] = 8'h00;
RAM[16'h7D5F] = 8'h00;
RAM[16'h7D60] = 8'h00;
RAM[16'h7D61] = 8'h00;
RAM[16'h7D62] = 8'h00;
RAM[16'h7D63] = 8'h00;
RAM[16'h7D64] = 8'h00;
RAM[16'h7D65] = 8'h00;
RAM[16'h7D66] = 8'h00;
RAM[16'h7D67] = 8'h00;
RAM[16'h7D68] = 8'h00;
RAM[16'h7D69] = 8'h00;
RAM[16'h7D6A] = 8'h00;
RAM[16'h7D6B] = 8'h00;
RAM[16'h7D6C] = 8'h00;
RAM[16'h7D6D] = 8'h00;
RAM[16'h7D6E] = 8'h00;
RAM[16'h7D6F] = 8'h00;
RAM[16'h7D70] = 8'h00;
RAM[16'h7D71] = 8'h00;
RAM[16'h7D72] = 8'h00;
RAM[16'h7D73] = 8'h00;
RAM[16'h7D74] = 8'h00;
RAM[16'h7D75] = 8'h00;
RAM[16'h7D76] = 8'h00;
RAM[16'h7D77] = 8'h00;
RAM[16'h7D78] = 8'h00;
RAM[16'h7D79] = 8'h00;
RAM[16'h7D7A] = 8'h00;
RAM[16'h7D7B] = 8'h00;
RAM[16'h7D7C] = 8'h00;
RAM[16'h7D7D] = 8'h00;
RAM[16'h7D7E] = 8'h00;
RAM[16'h7D7F] = 8'h00;
RAM[16'h7D80] = 8'h00;
RAM[16'h7D81] = 8'h00;
RAM[16'h7D82] = 8'h00;
RAM[16'h7D83] = 8'h00;
RAM[16'h7D84] = 8'h00;
RAM[16'h7D85] = 8'h00;
RAM[16'h7D86] = 8'h00;
RAM[16'h7D87] = 8'h00;
RAM[16'h7D88] = 8'h00;
RAM[16'h7D89] = 8'h00;
RAM[16'h7D8A] = 8'h00;
RAM[16'h7D8B] = 8'h00;
RAM[16'h7D8C] = 8'h00;
RAM[16'h7D8D] = 8'h00;
RAM[16'h7D8E] = 8'h00;
RAM[16'h7D8F] = 8'h00;
RAM[16'h7D90] = 8'h00;
RAM[16'h7D91] = 8'h00;
RAM[16'h7D92] = 8'h00;
RAM[16'h7D93] = 8'h00;
RAM[16'h7D94] = 8'h00;
RAM[16'h7D95] = 8'h00;
RAM[16'h7D96] = 8'h00;
RAM[16'h7D97] = 8'h00;
RAM[16'h7D98] = 8'h00;
RAM[16'h7D99] = 8'h00;
RAM[16'h7D9A] = 8'h00;
RAM[16'h7D9B] = 8'h00;
RAM[16'h7D9C] = 8'h00;
RAM[16'h7D9D] = 8'h00;
RAM[16'h7D9E] = 8'h00;
RAM[16'h7D9F] = 8'h00;
RAM[16'h7DA0] = 8'h00;
RAM[16'h7DA1] = 8'h00;
RAM[16'h7DA2] = 8'h00;
RAM[16'h7DA3] = 8'h00;
RAM[16'h7DA4] = 8'h00;
RAM[16'h7DA5] = 8'h00;
RAM[16'h7DA6] = 8'h00;
RAM[16'h7DA7] = 8'h00;
RAM[16'h7DA8] = 8'h00;
RAM[16'h7DA9] = 8'h00;
RAM[16'h7DAA] = 8'h00;
RAM[16'h7DAB] = 8'h00;
RAM[16'h7DAC] = 8'h00;
RAM[16'h7DAD] = 8'h00;
RAM[16'h7DAE] = 8'h00;
RAM[16'h7DAF] = 8'h00;
RAM[16'h7DB0] = 8'h00;
RAM[16'h7DB1] = 8'h00;
RAM[16'h7DB2] = 8'h00;
RAM[16'h7DB3] = 8'h00;
RAM[16'h7DB4] = 8'h00;
RAM[16'h7DB5] = 8'h00;
RAM[16'h7DB6] = 8'h00;
RAM[16'h7DB7] = 8'h00;
RAM[16'h7DB8] = 8'h00;
RAM[16'h7DB9] = 8'h00;
RAM[16'h7DBA] = 8'h00;
RAM[16'h7DBB] = 8'h00;
RAM[16'h7DBC] = 8'h00;
RAM[16'h7DBD] = 8'h00;
RAM[16'h7DBE] = 8'h00;
RAM[16'h7DBF] = 8'h00;
RAM[16'h7DC0] = 8'h00;
RAM[16'h7DC1] = 8'h00;
RAM[16'h7DC2] = 8'h00;
RAM[16'h7DC3] = 8'h00;
RAM[16'h7DC4] = 8'h00;
RAM[16'h7DC5] = 8'h00;
RAM[16'h7DC6] = 8'h00;
RAM[16'h7DC7] = 8'h00;
RAM[16'h7DC8] = 8'h00;
RAM[16'h7DC9] = 8'h00;
RAM[16'h7DCA] = 8'h00;
RAM[16'h7DCB] = 8'h00;
RAM[16'h7DCC] = 8'h00;
RAM[16'h7DCD] = 8'h00;
RAM[16'h7DCE] = 8'h00;
RAM[16'h7DCF] = 8'h00;
RAM[16'h7DD0] = 8'h00;
RAM[16'h7DD1] = 8'h00;
RAM[16'h7DD2] = 8'h00;
RAM[16'h7DD3] = 8'h00;
RAM[16'h7DD4] = 8'h00;
RAM[16'h7DD5] = 8'h00;
RAM[16'h7DD6] = 8'h00;
RAM[16'h7DD7] = 8'h00;
RAM[16'h7DD8] = 8'h00;
RAM[16'h7DD9] = 8'h00;
RAM[16'h7DDA] = 8'h00;
RAM[16'h7DDB] = 8'h00;
RAM[16'h7DDC] = 8'h00;
RAM[16'h7DDD] = 8'h00;
RAM[16'h7DDE] = 8'h00;
RAM[16'h7DDF] = 8'h00;
RAM[16'h7DE0] = 8'h00;
RAM[16'h7DE1] = 8'h00;
RAM[16'h7DE2] = 8'h00;
RAM[16'h7DE3] = 8'h00;
RAM[16'h7DE4] = 8'h00;
RAM[16'h7DE5] = 8'h00;
RAM[16'h7DE6] = 8'h00;
RAM[16'h7DE7] = 8'h00;
RAM[16'h7DE8] = 8'h00;
RAM[16'h7DE9] = 8'h00;
RAM[16'h7DEA] = 8'h00;
RAM[16'h7DEB] = 8'h00;
RAM[16'h7DEC] = 8'h00;
RAM[16'h7DED] = 8'h00;
RAM[16'h7DEE] = 8'h00;
RAM[16'h7DEF] = 8'h00;
RAM[16'h7DF0] = 8'h00;
RAM[16'h7DF1] = 8'h00;
RAM[16'h7DF2] = 8'h00;
RAM[16'h7DF3] = 8'h00;
RAM[16'h7DF4] = 8'h00;
RAM[16'h7DF5] = 8'h00;
RAM[16'h7DF6] = 8'h00;
RAM[16'h7DF7] = 8'h00;
RAM[16'h7DF8] = 8'h00;
RAM[16'h7DF9] = 8'h00;
RAM[16'h7DFA] = 8'h00;
RAM[16'h7DFB] = 8'h00;
RAM[16'h7DFC] = 8'h00;
RAM[16'h7DFD] = 8'h00;
RAM[16'h7DFE] = 8'h00;
RAM[16'h7DFF] = 8'h00;
RAM[16'h7E00] = 8'h00;
RAM[16'h7E01] = 8'h00;
RAM[16'h7E02] = 8'h00;
RAM[16'h7E03] = 8'h00;
RAM[16'h7E04] = 8'h00;
RAM[16'h7E05] = 8'h00;
RAM[16'h7E06] = 8'h00;
RAM[16'h7E07] = 8'h00;
RAM[16'h7E08] = 8'h00;
RAM[16'h7E09] = 8'h00;
RAM[16'h7E0A] = 8'h00;
RAM[16'h7E0B] = 8'h00;
RAM[16'h7E0C] = 8'h00;
RAM[16'h7E0D] = 8'h00;
RAM[16'h7E0E] = 8'h00;
RAM[16'h7E0F] = 8'h00;
RAM[16'h7E10] = 8'h00;
RAM[16'h7E11] = 8'h00;
RAM[16'h7E12] = 8'h00;
RAM[16'h7E13] = 8'h00;
RAM[16'h7E14] = 8'h00;
RAM[16'h7E15] = 8'h00;
RAM[16'h7E16] = 8'h00;
RAM[16'h7E17] = 8'h00;
RAM[16'h7E18] = 8'h00;
RAM[16'h7E19] = 8'h00;
RAM[16'h7E1A] = 8'h00;
RAM[16'h7E1B] = 8'h00;
RAM[16'h7E1C] = 8'h00;
RAM[16'h7E1D] = 8'h00;
RAM[16'h7E1E] = 8'h00;
RAM[16'h7E1F] = 8'h00;
RAM[16'h7E20] = 8'h00;
RAM[16'h7E21] = 8'h00;
RAM[16'h7E22] = 8'h00;
RAM[16'h7E23] = 8'h00;
RAM[16'h7E24] = 8'h00;
RAM[16'h7E25] = 8'h00;
RAM[16'h7E26] = 8'h00;
RAM[16'h7E27] = 8'h00;
RAM[16'h7E28] = 8'h00;
RAM[16'h7E29] = 8'h00;
RAM[16'h7E2A] = 8'h00;
RAM[16'h7E2B] = 8'h00;
RAM[16'h7E2C] = 8'h00;
RAM[16'h7E2D] = 8'h00;
RAM[16'h7E2E] = 8'h00;
RAM[16'h7E2F] = 8'h00;
RAM[16'h7E30] = 8'h00;
RAM[16'h7E31] = 8'h00;
RAM[16'h7E32] = 8'h00;
RAM[16'h7E33] = 8'h00;
RAM[16'h7E34] = 8'h00;
RAM[16'h7E35] = 8'h00;
RAM[16'h7E36] = 8'h00;
RAM[16'h7E37] = 8'h00;
RAM[16'h7E38] = 8'h00;
RAM[16'h7E39] = 8'h00;
RAM[16'h7E3A] = 8'h00;
RAM[16'h7E3B] = 8'h00;
RAM[16'h7E3C] = 8'h00;
RAM[16'h7E3D] = 8'h00;
RAM[16'h7E3E] = 8'h00;
RAM[16'h7E3F] = 8'h00;
RAM[16'h7E40] = 8'h00;
RAM[16'h7E41] = 8'h00;
RAM[16'h7E42] = 8'h00;
RAM[16'h7E43] = 8'h00;
RAM[16'h7E44] = 8'h00;
RAM[16'h7E45] = 8'h00;
RAM[16'h7E46] = 8'h00;
RAM[16'h7E47] = 8'h00;
RAM[16'h7E48] = 8'h00;
RAM[16'h7E49] = 8'h00;
RAM[16'h7E4A] = 8'h00;
RAM[16'h7E4B] = 8'h00;
RAM[16'h7E4C] = 8'h00;
RAM[16'h7E4D] = 8'h00;
RAM[16'h7E4E] = 8'h00;
RAM[16'h7E4F] = 8'h00;
RAM[16'h7E50] = 8'h00;
RAM[16'h7E51] = 8'h00;
RAM[16'h7E52] = 8'h00;
RAM[16'h7E53] = 8'h00;
RAM[16'h7E54] = 8'h00;
RAM[16'h7E55] = 8'h00;
RAM[16'h7E56] = 8'h00;
RAM[16'h7E57] = 8'h00;
RAM[16'h7E58] = 8'h00;
RAM[16'h7E59] = 8'h00;
RAM[16'h7E5A] = 8'h00;
RAM[16'h7E5B] = 8'h00;
RAM[16'h7E5C] = 8'h00;
RAM[16'h7E5D] = 8'h00;
RAM[16'h7E5E] = 8'h00;
RAM[16'h7E5F] = 8'h00;
RAM[16'h7E60] = 8'h00;
RAM[16'h7E61] = 8'h00;
RAM[16'h7E62] = 8'h00;
RAM[16'h7E63] = 8'h00;
RAM[16'h7E64] = 8'h00;
RAM[16'h7E65] = 8'h00;
RAM[16'h7E66] = 8'h00;
RAM[16'h7E67] = 8'h00;
RAM[16'h7E68] = 8'h00;
RAM[16'h7E69] = 8'h00;
RAM[16'h7E6A] = 8'h00;
RAM[16'h7E6B] = 8'h00;
RAM[16'h7E6C] = 8'h00;
RAM[16'h7E6D] = 8'h00;
RAM[16'h7E6E] = 8'h00;
RAM[16'h7E6F] = 8'h00;
RAM[16'h7E70] = 8'h00;
RAM[16'h7E71] = 8'h00;
RAM[16'h7E72] = 8'h00;
RAM[16'h7E73] = 8'h00;
RAM[16'h7E74] = 8'h00;
RAM[16'h7E75] = 8'h00;
RAM[16'h7E76] = 8'h00;
RAM[16'h7E77] = 8'h00;
RAM[16'h7E78] = 8'h00;
RAM[16'h7E79] = 8'h00;
RAM[16'h7E7A] = 8'h00;
RAM[16'h7E7B] = 8'h00;
RAM[16'h7E7C] = 8'h00;
RAM[16'h7E7D] = 8'h00;
RAM[16'h7E7E] = 8'h00;
RAM[16'h7E7F] = 8'h00;
RAM[16'h7E80] = 8'h00;
RAM[16'h7E81] = 8'h00;
RAM[16'h7E82] = 8'h00;
RAM[16'h7E83] = 8'h00;
RAM[16'h7E84] = 8'h00;
RAM[16'h7E85] = 8'h00;
RAM[16'h7E86] = 8'h00;
RAM[16'h7E87] = 8'h00;
RAM[16'h7E88] = 8'h00;
RAM[16'h7E89] = 8'h00;
RAM[16'h7E8A] = 8'h00;
RAM[16'h7E8B] = 8'h00;
RAM[16'h7E8C] = 8'h00;
RAM[16'h7E8D] = 8'h00;
RAM[16'h7E8E] = 8'h00;
RAM[16'h7E8F] = 8'h00;
RAM[16'h7E90] = 8'h00;
RAM[16'h7E91] = 8'h00;
RAM[16'h7E92] = 8'h00;
RAM[16'h7E93] = 8'h00;
RAM[16'h7E94] = 8'h00;
RAM[16'h7E95] = 8'h00;
RAM[16'h7E96] = 8'h00;
RAM[16'h7E97] = 8'h00;
RAM[16'h7E98] = 8'h00;
RAM[16'h7E99] = 8'h00;
RAM[16'h7E9A] = 8'h00;
RAM[16'h7E9B] = 8'h00;
RAM[16'h7E9C] = 8'h00;
RAM[16'h7E9D] = 8'h00;
RAM[16'h7E9E] = 8'h00;
RAM[16'h7E9F] = 8'h00;
RAM[16'h7EA0] = 8'h00;
RAM[16'h7EA1] = 8'h00;
RAM[16'h7EA2] = 8'h00;
RAM[16'h7EA3] = 8'h00;
RAM[16'h7EA4] = 8'h00;
RAM[16'h7EA5] = 8'h00;
RAM[16'h7EA6] = 8'h00;
RAM[16'h7EA7] = 8'h00;
RAM[16'h7EA8] = 8'h00;
RAM[16'h7EA9] = 8'h00;
RAM[16'h7EAA] = 8'h00;
RAM[16'h7EAB] = 8'h00;
RAM[16'h7EAC] = 8'h00;
RAM[16'h7EAD] = 8'h00;
RAM[16'h7EAE] = 8'h00;
RAM[16'h7EAF] = 8'h00;
RAM[16'h7EB0] = 8'h00;
RAM[16'h7EB1] = 8'h00;
RAM[16'h7EB2] = 8'h00;
RAM[16'h7EB3] = 8'h00;
RAM[16'h7EB4] = 8'h00;
RAM[16'h7EB5] = 8'h00;
RAM[16'h7EB6] = 8'h00;
RAM[16'h7EB7] = 8'h00;
RAM[16'h7EB8] = 8'h00;
RAM[16'h7EB9] = 8'h00;
RAM[16'h7EBA] = 8'h00;
RAM[16'h7EBB] = 8'h00;
RAM[16'h7EBC] = 8'h00;
RAM[16'h7EBD] = 8'h00;
RAM[16'h7EBE] = 8'h00;
RAM[16'h7EBF] = 8'h00;
RAM[16'h7EC0] = 8'h00;
RAM[16'h7EC1] = 8'h00;
RAM[16'h7EC2] = 8'h00;
RAM[16'h7EC3] = 8'h00;
RAM[16'h7EC4] = 8'h00;
RAM[16'h7EC5] = 8'h00;
RAM[16'h7EC6] = 8'h00;
RAM[16'h7EC7] = 8'h00;
RAM[16'h7EC8] = 8'h00;
RAM[16'h7EC9] = 8'h00;
RAM[16'h7ECA] = 8'h00;
RAM[16'h7ECB] = 8'h00;
RAM[16'h7ECC] = 8'h00;
RAM[16'h7ECD] = 8'h00;
RAM[16'h7ECE] = 8'h00;
RAM[16'h7ECF] = 8'h00;
RAM[16'h7ED0] = 8'h00;
RAM[16'h7ED1] = 8'h00;
RAM[16'h7ED2] = 8'h00;
RAM[16'h7ED3] = 8'h00;
RAM[16'h7ED4] = 8'h00;
RAM[16'h7ED5] = 8'h00;
RAM[16'h7ED6] = 8'h00;
RAM[16'h7ED7] = 8'h00;
RAM[16'h7ED8] = 8'h00;
RAM[16'h7ED9] = 8'h00;
RAM[16'h7EDA] = 8'h00;
RAM[16'h7EDB] = 8'h00;
RAM[16'h7EDC] = 8'h00;
RAM[16'h7EDD] = 8'h00;
RAM[16'h7EDE] = 8'h00;
RAM[16'h7EDF] = 8'h00;
RAM[16'h7EE0] = 8'h00;
RAM[16'h7EE1] = 8'h00;
RAM[16'h7EE2] = 8'h00;
RAM[16'h7EE3] = 8'h00;
RAM[16'h7EE4] = 8'h00;
RAM[16'h7EE5] = 8'h00;
RAM[16'h7EE6] = 8'h00;
RAM[16'h7EE7] = 8'h00;
RAM[16'h7EE8] = 8'h00;
RAM[16'h7EE9] = 8'h00;
RAM[16'h7EEA] = 8'h00;
RAM[16'h7EEB] = 8'h00;
RAM[16'h7EEC] = 8'h00;
RAM[16'h7EED] = 8'h00;
RAM[16'h7EEE] = 8'h00;
RAM[16'h7EEF] = 8'h00;
RAM[16'h7EF0] = 8'h00;
RAM[16'h7EF1] = 8'h00;
RAM[16'h7EF2] = 8'h00;
RAM[16'h7EF3] = 8'h00;
RAM[16'h7EF4] = 8'h00;
RAM[16'h7EF5] = 8'h00;
RAM[16'h7EF6] = 8'h00;
RAM[16'h7EF7] = 8'h00;
RAM[16'h7EF8] = 8'h00;
RAM[16'h7EF9] = 8'h00;
RAM[16'h7EFA] = 8'h00;
RAM[16'h7EFB] = 8'h00;
RAM[16'h7EFC] = 8'h00;
RAM[16'h7EFD] = 8'h00;
RAM[16'h7EFE] = 8'h00;
RAM[16'h7EFF] = 8'h00;
RAM[16'h7F00] = 8'h00;
RAM[16'h7F01] = 8'h00;
RAM[16'h7F02] = 8'h00;
RAM[16'h7F03] = 8'h00;
RAM[16'h7F04] = 8'h00;
RAM[16'h7F05] = 8'h00;
RAM[16'h7F06] = 8'h00;
RAM[16'h7F07] = 8'h00;
RAM[16'h7F08] = 8'h00;
RAM[16'h7F09] = 8'h00;
RAM[16'h7F0A] = 8'h00;
RAM[16'h7F0B] = 8'h00;
RAM[16'h7F0C] = 8'h00;
RAM[16'h7F0D] = 8'h00;
RAM[16'h7F0E] = 8'h00;
RAM[16'h7F0F] = 8'h00;
RAM[16'h7F10] = 8'h00;
RAM[16'h7F11] = 8'h00;
RAM[16'h7F12] = 8'h00;
RAM[16'h7F13] = 8'h00;
RAM[16'h7F14] = 8'h00;
RAM[16'h7F15] = 8'h00;
RAM[16'h7F16] = 8'h00;
RAM[16'h7F17] = 8'h00;
RAM[16'h7F18] = 8'h00;
RAM[16'h7F19] = 8'h00;
RAM[16'h7F1A] = 8'h00;
RAM[16'h7F1B] = 8'h00;
RAM[16'h7F1C] = 8'h00;
RAM[16'h7F1D] = 8'h00;
RAM[16'h7F1E] = 8'h00;
RAM[16'h7F1F] = 8'h00;
RAM[16'h7F20] = 8'h00;
RAM[16'h7F21] = 8'h00;
RAM[16'h7F22] = 8'h00;
RAM[16'h7F23] = 8'h00;
RAM[16'h7F24] = 8'h00;
RAM[16'h7F25] = 8'h00;
RAM[16'h7F26] = 8'h00;
RAM[16'h7F27] = 8'h00;
RAM[16'h7F28] = 8'h00;
RAM[16'h7F29] = 8'h00;
RAM[16'h7F2A] = 8'h00;
RAM[16'h7F2B] = 8'h00;
RAM[16'h7F2C] = 8'h00;
RAM[16'h7F2D] = 8'h00;
RAM[16'h7F2E] = 8'h00;
RAM[16'h7F2F] = 8'h00;
RAM[16'h7F30] = 8'h00;
RAM[16'h7F31] = 8'h00;
RAM[16'h7F32] = 8'h00;
RAM[16'h7F33] = 8'h00;
RAM[16'h7F34] = 8'h00;
RAM[16'h7F35] = 8'h00;
RAM[16'h7F36] = 8'h00;
RAM[16'h7F37] = 8'h00;
RAM[16'h7F38] = 8'h00;
RAM[16'h7F39] = 8'h00;
RAM[16'h7F3A] = 8'h00;
RAM[16'h7F3B] = 8'h00;
RAM[16'h7F3C] = 8'h00;
RAM[16'h7F3D] = 8'h00;
RAM[16'h7F3E] = 8'h00;
RAM[16'h7F3F] = 8'h00;
RAM[16'h7F40] = 8'h00;
RAM[16'h7F41] = 8'h00;
RAM[16'h7F42] = 8'h00;
RAM[16'h7F43] = 8'h00;
RAM[16'h7F44] = 8'h00;
RAM[16'h7F45] = 8'h00;
RAM[16'h7F46] = 8'h00;
RAM[16'h7F47] = 8'h00;
RAM[16'h7F48] = 8'h00;
RAM[16'h7F49] = 8'h00;
RAM[16'h7F4A] = 8'h00;
RAM[16'h7F4B] = 8'h00;
RAM[16'h7F4C] = 8'h00;
RAM[16'h7F4D] = 8'h00;
RAM[16'h7F4E] = 8'h00;
RAM[16'h7F4F] = 8'h00;
RAM[16'h7F50] = 8'h00;
RAM[16'h7F51] = 8'h00;
RAM[16'h7F52] = 8'h00;
RAM[16'h7F53] = 8'h00;
RAM[16'h7F54] = 8'h00;
RAM[16'h7F55] = 8'h00;
RAM[16'h7F56] = 8'h00;
RAM[16'h7F57] = 8'h00;
RAM[16'h7F58] = 8'h00;
RAM[16'h7F59] = 8'h00;
RAM[16'h7F5A] = 8'h00;
RAM[16'h7F5B] = 8'h00;
RAM[16'h7F5C] = 8'h00;
RAM[16'h7F5D] = 8'h00;
RAM[16'h7F5E] = 8'h00;
RAM[16'h7F5F] = 8'h00;
RAM[16'h7F60] = 8'h00;
RAM[16'h7F61] = 8'h00;
RAM[16'h7F62] = 8'h00;
RAM[16'h7F63] = 8'h00;
RAM[16'h7F64] = 8'h00;
RAM[16'h7F65] = 8'h00;
RAM[16'h7F66] = 8'h00;
RAM[16'h7F67] = 8'h00;
RAM[16'h7F68] = 8'h00;
RAM[16'h7F69] = 8'h00;
RAM[16'h7F6A] = 8'h00;
RAM[16'h7F6B] = 8'h00;
RAM[16'h7F6C] = 8'h00;
RAM[16'h7F6D] = 8'h00;
RAM[16'h7F6E] = 8'h00;
RAM[16'h7F6F] = 8'h00;
RAM[16'h7F70] = 8'h00;
RAM[16'h7F71] = 8'h00;
RAM[16'h7F72] = 8'h00;
RAM[16'h7F73] = 8'h00;
RAM[16'h7F74] = 8'h00;
RAM[16'h7F75] = 8'h00;
RAM[16'h7F76] = 8'h00;
RAM[16'h7F77] = 8'h00;
RAM[16'h7F78] = 8'h00;
RAM[16'h7F79] = 8'h00;
RAM[16'h7F7A] = 8'h00;
RAM[16'h7F7B] = 8'h00;
RAM[16'h7F7C] = 8'h00;
RAM[16'h7F7D] = 8'h00;
RAM[16'h7F7E] = 8'h00;
RAM[16'h7F7F] = 8'h00;
RAM[16'h7F80] = 8'h00;
RAM[16'h7F81] = 8'h00;
RAM[16'h7F82] = 8'h00;
RAM[16'h7F83] = 8'h00;
RAM[16'h7F84] = 8'h00;
RAM[16'h7F85] = 8'h00;
RAM[16'h7F86] = 8'h00;
RAM[16'h7F87] = 8'h00;
RAM[16'h7F88] = 8'h00;
RAM[16'h7F89] = 8'h00;
RAM[16'h7F8A] = 8'h00;
RAM[16'h7F8B] = 8'h00;
RAM[16'h7F8C] = 8'h00;
RAM[16'h7F8D] = 8'h00;
RAM[16'h7F8E] = 8'h00;
RAM[16'h7F8F] = 8'h00;
RAM[16'h7F90] = 8'h00;
RAM[16'h7F91] = 8'h00;
RAM[16'h7F92] = 8'h00;
RAM[16'h7F93] = 8'h00;
RAM[16'h7F94] = 8'h00;
RAM[16'h7F95] = 8'h00;
RAM[16'h7F96] = 8'h00;
RAM[16'h7F97] = 8'h00;
RAM[16'h7F98] = 8'h00;
RAM[16'h7F99] = 8'h00;
RAM[16'h7F9A] = 8'h00;
RAM[16'h7F9B] = 8'h00;
RAM[16'h7F9C] = 8'h00;
RAM[16'h7F9D] = 8'h00;
RAM[16'h7F9E] = 8'h00;
RAM[16'h7F9F] = 8'h00;
RAM[16'h7FA0] = 8'h00;
RAM[16'h7FA1] = 8'h00;
RAM[16'h7FA2] = 8'h00;
RAM[16'h7FA3] = 8'h00;
RAM[16'h7FA4] = 8'h00;
RAM[16'h7FA5] = 8'h00;
RAM[16'h7FA6] = 8'h00;
RAM[16'h7FA7] = 8'h00;
RAM[16'h7FA8] = 8'h00;
RAM[16'h7FA9] = 8'h00;
RAM[16'h7FAA] = 8'h00;
RAM[16'h7FAB] = 8'h00;
RAM[16'h7FAC] = 8'h00;
RAM[16'h7FAD] = 8'h00;
RAM[16'h7FAE] = 8'h00;
RAM[16'h7FAF] = 8'h00;
RAM[16'h7FB0] = 8'h00;
RAM[16'h7FB1] = 8'h00;
RAM[16'h7FB2] = 8'h00;
RAM[16'h7FB3] = 8'h00;
RAM[16'h7FB4] = 8'h00;
RAM[16'h7FB5] = 8'h00;
RAM[16'h7FB6] = 8'h00;
RAM[16'h7FB7] = 8'h00;
RAM[16'h7FB8] = 8'h00;
RAM[16'h7FB9] = 8'h00;
RAM[16'h7FBA] = 8'h00;
RAM[16'h7FBB] = 8'h00;
RAM[16'h7FBC] = 8'h00;
RAM[16'h7FBD] = 8'h00;
RAM[16'h7FBE] = 8'h00;
RAM[16'h7FBF] = 8'h00;
RAM[16'h7FC0] = 8'h00;
RAM[16'h7FC1] = 8'h00;
RAM[16'h7FC2] = 8'h00;
RAM[16'h7FC3] = 8'h00;
RAM[16'h7FC4] = 8'h00;
RAM[16'h7FC5] = 8'h00;
RAM[16'h7FC6] = 8'h00;
RAM[16'h7FC7] = 8'h00;
RAM[16'h7FC8] = 8'h00;
RAM[16'h7FC9] = 8'h00;
RAM[16'h7FCA] = 8'h00;
RAM[16'h7FCB] = 8'h00;
RAM[16'h7FCC] = 8'h00;
RAM[16'h7FCD] = 8'h00;
RAM[16'h7FCE] = 8'h00;
RAM[16'h7FCF] = 8'h00;
RAM[16'h7FD0] = 8'h00;
RAM[16'h7FD1] = 8'h00;
RAM[16'h7FD2] = 8'h00;
RAM[16'h7FD3] = 8'h00;
RAM[16'h7FD4] = 8'h00;
RAM[16'h7FD5] = 8'h00;
RAM[16'h7FD6] = 8'h00;
RAM[16'h7FD7] = 8'h00;
RAM[16'h7FD8] = 8'h00;
RAM[16'h7FD9] = 8'h00;
RAM[16'h7FDA] = 8'h00;
RAM[16'h7FDB] = 8'h00;
RAM[16'h7FDC] = 8'h00;
RAM[16'h7FDD] = 8'h00;
RAM[16'h7FDE] = 8'h00;
RAM[16'h7FDF] = 8'h00;
RAM[16'h7FE0] = 8'h00;
RAM[16'h7FE1] = 8'h00;
RAM[16'h7FE2] = 8'h00;
RAM[16'h7FE3] = 8'h00;
RAM[16'h7FE4] = 8'h00;
RAM[16'h7FE5] = 8'h00;
RAM[16'h7FE6] = 8'h00;
RAM[16'h7FE7] = 8'h00;
RAM[16'h7FE8] = 8'h00;
RAM[16'h7FE9] = 8'h00;
RAM[16'h7FEA] = 8'h00;
RAM[16'h7FEB] = 8'h00;
RAM[16'h7FEC] = 8'h00;
RAM[16'h7FED] = 8'h00;
RAM[16'h7FEE] = 8'h00;
RAM[16'h7FEF] = 8'h00;
RAM[16'h7FF0] = 8'h00;
RAM[16'h7FF1] = 8'h00;
RAM[16'h7FF2] = 8'h00;
RAM[16'h7FF3] = 8'h00;
RAM[16'h7FF4] = 8'h00;
RAM[16'h7FF5] = 8'h00;
RAM[16'h7FF6] = 8'h00;
RAM[16'h7FF7] = 8'h00;
RAM[16'h7FF8] = 8'h00;
RAM[16'h7FF9] = 8'h00;
RAM[16'h7FFA] = 8'h00;
RAM[16'h7FFB] = 8'h00;
RAM[16'h7FFC] = 8'h00;
RAM[16'h7FFD] = 8'h00;
RAM[16'h7FFE] = 8'h00;
RAM[16'h7FFF] = 8'h00;
end
