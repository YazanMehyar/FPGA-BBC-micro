`define KiB16 16383
`define KiB32 32767
`define KiB64 65535
`define CLKPERIOD 10

`timescale 1ns/1ns
