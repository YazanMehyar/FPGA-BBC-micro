initial begin
DFS[16'h0000] = 8'h00;
DFS[16'h0001] = 8'h00;
DFS[16'h0002] = 8'h00;
DFS[16'h0003] = 8'h4C;
DFS[16'h0004] = 8'h55;
DFS[16'h0005] = 8'h94;
DFS[16'h0006] = 8'h82;
DFS[16'h0007] = 8'h11;
DFS[16'h0008] = 8'h5A;
DFS[16'h0009] = 8'h44;
DFS[16'h000A] = 8'h46;
DFS[16'h000B] = 8'h53;
DFS[16'h000C] = 8'h00;
DFS[16'h000D] = 8'h30;
DFS[16'h000E] = 8'h2E;
DFS[16'h000F] = 8'h39;
DFS[16'h0010] = 8'h30;
DFS[16'h0011] = 8'h00;
DFS[16'h0012] = 8'h28;
DFS[16'h0013] = 8'h43;
DFS[16'h0014] = 8'h29;
DFS[16'h0015] = 8'h6C;
DFS[16'h0016] = 8'h1E;
DFS[16'h0017] = 8'h02;
DFS[16'h0018] = 8'h20;
DFS[16'h0019] = 8'h5B;
DFS[16'h001A] = 8'h80;
DFS[16'h001B] = 8'h44;
DFS[16'h001C] = 8'h69;
DFS[16'h001D] = 8'h73;
DFS[16'h001E] = 8'h6B;
DFS[16'h001F] = 8'h20;
DFS[16'h0020] = 8'h90;
DFS[16'h0021] = 8'h11;
DFS[16'h0022] = 8'h20;
DFS[16'h0023] = 8'h5B;
DFS[16'h0024] = 8'h80;
DFS[16'h0025] = 8'h42;
DFS[16'h0026] = 8'h61;
DFS[16'h0027] = 8'h64;
DFS[16'h0028] = 8'h20;
DFS[16'h0029] = 8'h90;
DFS[16'h002A] = 8'h08;
DFS[16'h002B] = 8'h20;
DFS[16'h002C] = 8'h5B;
DFS[16'h002D] = 8'h80;
DFS[16'h002E] = 8'h46;
DFS[16'h002F] = 8'h69;
DFS[16'h0030] = 8'h6C;
DFS[16'h0031] = 8'h65;
DFS[16'h0032] = 8'h20;
DFS[16'h0033] = 8'h85;
DFS[16'h0034] = 8'hB3;
DFS[16'h0035] = 8'h68;
DFS[16'h0036] = 8'h85;
DFS[16'h0037] = 8'hAE;
DFS[16'h0038] = 8'h68;
DFS[16'h0039] = 8'h85;
DFS[16'h003A] = 8'hAF;
DFS[16'h003B] = 8'hA5;
DFS[16'h003C] = 8'hB3;
DFS[16'h003D] = 8'h48;
DFS[16'h003E] = 8'h98;
DFS[16'h003F] = 8'h48;
DFS[16'h0040] = 8'hA0;
DFS[16'h0041] = 8'h00;
DFS[16'h0042] = 8'h20;
DFS[16'h0043] = 8'hDA;
DFS[16'h0044] = 8'h83;
DFS[16'h0045] = 8'hB1;
DFS[16'h0046] = 8'hAE;
DFS[16'h0047] = 8'h8D;
DFS[16'h0048] = 8'h01;
DFS[16'h0049] = 8'h01;
DFS[16'h004A] = 8'h2C;
DFS[16'h004B] = 8'hDE;
DFS[16'h004C] = 8'h10;
DFS[16'h004D] = 8'h10;
DFS[16'h004E] = 8'h25;
DFS[16'h004F] = 8'hA9;
DFS[16'h0050] = 8'h02;
DFS[16'h0051] = 8'h8D;
DFS[16'h0052] = 8'hDE;
DFS[16'h0053] = 8'h10;
DFS[16'h0054] = 8'hA9;
DFS[16'h0055] = 8'h00;
DFS[16'h0056] = 8'h8D;
DFS[16'h0057] = 8'h00;
DFS[16'h0058] = 8'h01;
DFS[16'h0059] = 8'hF0;
DFS[16'h005A] = 8'h19;
DFS[16'h005B] = 8'hA9;
DFS[16'h005C] = 8'h02;
DFS[16'h005D] = 8'h8D;
DFS[16'h005E] = 8'hDE;
DFS[16'h005F] = 8'h10;
DFS[16'h0060] = 8'hA9;
DFS[16'h0061] = 8'h00;
DFS[16'h0062] = 8'h8D;
DFS[16'h0063] = 8'h00;
DFS[16'h0064] = 8'h01;
DFS[16'h0065] = 8'h85;
DFS[16'h0066] = 8'hB3;
DFS[16'h0067] = 8'h68;
DFS[16'h0068] = 8'h85;
DFS[16'h0069] = 8'hAE;
DFS[16'h006A] = 8'h68;
DFS[16'h006B] = 8'h85;
DFS[16'h006C] = 8'hAF;
DFS[16'h006D] = 8'hA5;
DFS[16'h006E] = 8'hB3;
DFS[16'h006F] = 8'h48;
DFS[16'h0070] = 8'h98;
DFS[16'h0071] = 8'h48;
DFS[16'h0072] = 8'hA0;
DFS[16'h0073] = 8'h00;
DFS[16'h0074] = 8'h20;
DFS[16'h0075] = 8'hDA;
DFS[16'h0076] = 8'h83;
DFS[16'h0077] = 8'hB1;
DFS[16'h0078] = 8'hAE;
DFS[16'h0079] = 8'h30;
DFS[16'h007A] = 8'h08;
DFS[16'h007B] = 8'hF0;
DFS[16'h007C] = 8'h0D;
DFS[16'h007D] = 8'h20;
DFS[16'h007E] = 8'h9C;
DFS[16'h007F] = 8'h80;
DFS[16'h0080] = 8'h4C;
DFS[16'h0081] = 8'h74;
DFS[16'h0082] = 8'h80;
DFS[16'h0083] = 8'h68;
DFS[16'h0084] = 8'hA8;
DFS[16'h0085] = 8'h68;
DFS[16'h0086] = 8'h18;
DFS[16'h0087] = 8'h6C;
DFS[16'h0088] = 8'hAE;
DFS[16'h0089] = 8'h00;
DFS[16'h008A] = 8'hA9;
DFS[16'h008B] = 8'h00;
DFS[16'h008C] = 8'hAE;
DFS[16'h008D] = 8'hDE;
DFS[16'h008E] = 8'h10;
DFS[16'h008F] = 8'h9D;
DFS[16'h0090] = 8'h00;
DFS[16'h0091] = 8'h01;
DFS[16'h0092] = 8'hA9;
DFS[16'h0093] = 8'hFF;
DFS[16'h0094] = 8'h8D;
DFS[16'h0095] = 8'hDE;
DFS[16'h0096] = 8'h10;
DFS[16'h0097] = 8'h4C;
DFS[16'h0098] = 8'h00;
DFS[16'h0099] = 8'h01;
DFS[16'h009A] = 8'hA9;
DFS[16'h009B] = 8'h2E;
DFS[16'h009C] = 8'h20;
DFS[16'h009D] = 8'hE1;
DFS[16'h009E] = 8'h83;
DFS[16'h009F] = 8'h2C;
DFS[16'h00A0] = 8'hDE;
DFS[16'h00A1] = 8'h10;
DFS[16'h00A2] = 8'h10;
DFS[16'h00A3] = 8'h14;
DFS[16'h00A4] = 8'h48;
DFS[16'h00A5] = 8'h20;
DFS[16'h00A6] = 8'h1C;
DFS[16'h00A7] = 8'h99;
DFS[16'h00A8] = 8'h8A;
DFS[16'h00A9] = 8'h48;
DFS[16'h00AA] = 8'h09;
DFS[16'h00AB] = 8'h10;
DFS[16'h00AC] = 8'h20;
DFS[16'h00AD] = 8'h17;
DFS[16'h00AE] = 8'h99;
DFS[16'h00AF] = 8'h68;
DFS[16'h00B0] = 8'hAA;
DFS[16'h00B1] = 8'h68;
DFS[16'h00B2] = 8'h20;
DFS[16'h00B3] = 8'hE3;
DFS[16'h00B4] = 8'hFF;
DFS[16'h00B5] = 8'h4C;
DFS[16'h00B6] = 8'h18;
DFS[16'h00B7] = 8'h99;
DFS[16'h00B8] = 8'hAE;
DFS[16'h00B9] = 8'hDE;
DFS[16'h00BA] = 8'h10;
DFS[16'h00BB] = 8'h9D;
DFS[16'h00BC] = 8'h00;
DFS[16'h00BD] = 8'h01;
DFS[16'h00BE] = 8'hEE;
DFS[16'h00BF] = 8'hDE;
DFS[16'h00C0] = 8'h10;
DFS[16'h00C1] = 8'h60;
DFS[16'h00C2] = 8'h48;
DFS[16'h00C3] = 8'h20;
DFS[16'h00C4] = 8'h05;
DFS[16'h00C5] = 8'h82;
DFS[16'h00C6] = 8'h20;
DFS[16'h00C7] = 8'hCA;
DFS[16'h00C8] = 8'h80;
DFS[16'h00C9] = 8'h68;
DFS[16'h00CA] = 8'h48;
DFS[16'h00CB] = 8'h29;
DFS[16'h00CC] = 8'h0F;
DFS[16'h00CD] = 8'hC9;
DFS[16'h00CE] = 8'h0A;
DFS[16'h00CF] = 8'h90;
DFS[16'h00D0] = 8'h02;
DFS[16'h00D1] = 8'h69;
DFS[16'h00D2] = 8'h06;
DFS[16'h00D3] = 8'h69;
DFS[16'h00D4] = 8'h30;
DFS[16'h00D5] = 8'h20;
DFS[16'h00D6] = 8'h9C;
DFS[16'h00D7] = 8'h80;
DFS[16'h00D8] = 8'h68;
DFS[16'h00D9] = 8'h60;
DFS[16'h00DA] = 8'h20;
DFS[16'h00DB] = 8'hEA;
DFS[16'h00DC] = 8'h80;
DFS[16'h00DD] = 8'hCA;
DFS[16'h00DE] = 8'hCA;
DFS[16'h00DF] = 8'h20;
DFS[16'h00E0] = 8'hE2;
DFS[16'h00E1] = 8'h80;
DFS[16'h00E2] = 8'hB1;
DFS[16'h00E3] = 8'hB0;
DFS[16'h00E4] = 8'h9D;
DFS[16'h00E5] = 8'h72;
DFS[16'h00E6] = 8'h10;
DFS[16'h00E7] = 8'hE8;
DFS[16'h00E8] = 8'hC8;
DFS[16'h00E9] = 8'h60;
DFS[16'h00EA] = 8'h20;
DFS[16'h00EB] = 8'hED;
DFS[16'h00EC] = 8'h80;
DFS[16'h00ED] = 8'hB1;
DFS[16'h00EE] = 8'hB0;
DFS[16'h00EF] = 8'h95;
DFS[16'h00F0] = 8'hBC;
DFS[16'h00F1] = 8'hE8;
DFS[16'h00F2] = 8'hC8;
DFS[16'h00F3] = 8'h60;
DFS[16'h00F4] = 8'hA9;
DFS[16'h00F5] = 8'h20;
DFS[16'h00F6] = 8'hA2;
DFS[16'h00F7] = 8'h06;
DFS[16'h00F8] = 8'h95;
DFS[16'h00F9] = 8'hC7;
DFS[16'h00FA] = 8'hCA;
DFS[16'h00FB] = 8'h10;
DFS[16'h00FC] = 8'hFB;
DFS[16'h00FD] = 8'h60;
DFS[16'h00FE] = 8'h20;
DFS[16'h00FF] = 8'h4D;
DFS[16'h0100] = 8'h83;
DFS[16'h0101] = 8'h20;
DFS[16'h0102] = 8'hF4;
DFS[16'h0103] = 8'h80;
DFS[16'h0104] = 8'h30;
DFS[16'h0105] = 8'h13;
DFS[16'h0106] = 8'h20;
DFS[16'h0107] = 8'h4D;
DFS[16'h0108] = 8'h83;
DFS[16'h0109] = 8'h20;
DFS[16'h010A] = 8'hF4;
DFS[16'h010B] = 8'h80;
DFS[16'h010C] = 8'hA5;
DFS[16'h010D] = 8'hBC;
DFS[16'h010E] = 8'h85;
DFS[16'h010F] = 8'hF2;
DFS[16'h0110] = 8'hA5;
DFS[16'h0111] = 8'hBD;
DFS[16'h0112] = 8'h85;
DFS[16'h0113] = 8'hF3;
DFS[16'h0114] = 8'hA0;
DFS[16'h0115] = 8'h00;
DFS[16'h0116] = 8'h20;
DFS[16'h0117] = 8'hBF;
DFS[16'h0118] = 8'h86;
DFS[16'h0119] = 8'hA2;
DFS[16'h011A] = 8'h01;
DFS[16'h011B] = 8'h20;
DFS[16'h011C] = 8'hC5;
DFS[16'h011D] = 8'hFF;
DFS[16'h011E] = 8'hB0;
DFS[16'h011F] = 8'hDD;
DFS[16'h0120] = 8'h85;
DFS[16'h0121] = 8'hC7;
DFS[16'h0122] = 8'hC9;
DFS[16'h0123] = 8'h2E;
DFS[16'h0124] = 8'hD0;
DFS[16'h0125] = 8'h04;
DFS[16'h0126] = 8'hA9;
DFS[16'h0127] = 8'h20;
DFS[16'h0128] = 8'hD0;
DFS[16'h0129] = 8'h4D;
DFS[16'h012A] = 8'hC9;
DFS[16'h012B] = 8'h3A;
DFS[16'h012C] = 8'hD0;
DFS[16'h012D] = 8'h21;
DFS[16'h012E] = 8'h20;
DFS[16'h012F] = 8'hC5;
DFS[16'h0130] = 8'hFF;
DFS[16'h0131] = 8'hB0;
DFS[16'h0132] = 8'h15;
DFS[16'h0133] = 8'h38;
DFS[16'h0134] = 8'hE9;
DFS[16'h0135] = 8'h30;
DFS[16'h0136] = 8'h90;
DFS[16'h0137] = 8'h10;
DFS[16'h0138] = 8'hC9;
DFS[16'h0139] = 8'h04;
DFS[16'h013A] = 8'hB0;
DFS[16'h013B] = 8'h0C;
DFS[16'h013C] = 8'h20;
DFS[16'h013D] = 8'h7E;
DFS[16'h013E] = 8'h87;
DFS[16'h013F] = 8'h20;
DFS[16'h0140] = 8'hC5;
DFS[16'h0141] = 8'hFF;
DFS[16'h0142] = 8'hB0;
DFS[16'h0143] = 8'h5C;
DFS[16'h0144] = 8'hC9;
DFS[16'h0145] = 8'h2E;
DFS[16'h0146] = 8'hF0;
DFS[16'h0147] = 8'h03;
DFS[16'h0148] = 8'h4C;
DFS[16'h0149] = 8'h74;
DFS[16'h014A] = 8'h83;
DFS[16'h014B] = 8'hA9;
DFS[16'h014C] = 8'h24;
DFS[16'h014D] = 8'hD0;
DFS[16'h014E] = 8'h28;
DFS[16'h014F] = 8'hC9;
DFS[16'h0150] = 8'h2A;
DFS[16'h0151] = 8'hD0;
DFS[16'h0152] = 8'h19;
DFS[16'h0153] = 8'h20;
DFS[16'h0154] = 8'hC5;
DFS[16'h0155] = 8'hFF;
DFS[16'h0156] = 8'hB0;
DFS[16'h0157] = 8'h08;
DFS[16'h0158] = 8'hC9;
DFS[16'h0159] = 8'h2E;
DFS[16'h015A] = 8'hD0;
DFS[16'h015B] = 8'h32;
DFS[16'h015C] = 8'hA9;
DFS[16'h015D] = 8'h23;
DFS[16'h015E] = 8'hD0;
DFS[16'h015F] = 8'h17;
DFS[16'h0160] = 8'hA2;
DFS[16'h0161] = 8'h00;
DFS[16'h0162] = 8'hA9;
DFS[16'h0163] = 8'h23;
DFS[16'h0164] = 8'h95;
DFS[16'h0165] = 8'hC7;
DFS[16'h0166] = 8'hE8;
DFS[16'h0167] = 8'hE0;
DFS[16'h0168] = 8'h07;
DFS[16'h0169] = 8'hD0;
DFS[16'h016A] = 8'hF9;
DFS[16'h016B] = 8'h60;
DFS[16'h016C] = 8'h20;
DFS[16'h016D] = 8'hC5;
DFS[16'h016E] = 8'hFF;
DFS[16'h016F] = 8'hB0;
DFS[16'h0170] = 8'h2F;
DFS[16'h0171] = 8'hC9;
DFS[16'h0172] = 8'h2E;
DFS[16'h0173] = 8'hD0;
DFS[16'h0174] = 8'h10;
DFS[16'h0175] = 8'hA5;
DFS[16'h0176] = 8'hC7;
DFS[16'h0177] = 8'h85;
DFS[16'h0178] = 8'hCE;
DFS[16'h0179] = 8'h4C;
DFS[16'h017A] = 8'h1B;
DFS[16'h017B] = 8'h81;
DFS[16'h017C] = 8'h20;
DFS[16'h017D] = 8'hC5;
DFS[16'h017E] = 8'hFF;
DFS[16'h017F] = 8'hB0;
DFS[16'h0180] = 8'h1F;
DFS[16'h0181] = 8'hE0;
DFS[16'h0182] = 8'h07;
DFS[16'h0183] = 8'hF0;
DFS[16'h0184] = 8'h09;
DFS[16'h0185] = 8'hC9;
DFS[16'h0186] = 8'h2A;
DFS[16'h0187] = 8'hD0;
DFS[16'h0188] = 8'h12;
DFS[16'h0189] = 8'h20;
DFS[16'h018A] = 8'hC5;
DFS[16'h018B] = 8'hFF;
DFS[16'h018C] = 8'hB0;
DFS[16'h018D] = 8'hD4;
DFS[16'h018E] = 8'h20;
DFS[16'h018F] = 8'h22;
DFS[16'h0190] = 8'h80;
DFS[16'h0191] = 8'hCC;
DFS[16'h0192] = 8'h66;
DFS[16'h0193] = 8'h69;
DFS[16'h0194] = 8'h6C;
DFS[16'h0195] = 8'h65;
DFS[16'h0196] = 8'h6E;
DFS[16'h0197] = 8'h61;
DFS[16'h0198] = 8'h6D;
DFS[16'h0199] = 8'h65;
DFS[16'h019A] = 8'h00;
DFS[16'h019B] = 8'h95;
DFS[16'h019C] = 8'hC7;
DFS[16'h019D] = 8'hE8;
DFS[16'h019E] = 8'hD0;
DFS[16'h019F] = 8'hDC;
DFS[16'h01A0] = 8'h60;
DFS[16'h01A1] = 8'h20;
DFS[16'h01A2] = 8'hE1;
DFS[16'h01A3] = 8'h83;
DFS[16'h01A4] = 8'hAD;
DFS[16'h01A5] = 8'h04;
DFS[16'h01A6] = 8'h0F;
DFS[16'h01A7] = 8'h20;
DFS[16'h01A8] = 8'h47;
DFS[16'h01A9] = 8'h83;
DFS[16'h01AA] = 8'hCD;
DFS[16'h01AB] = 8'h04;
DFS[16'h01AC] = 8'h0F;
DFS[16'h01AD] = 8'hF0;
DFS[16'h01AE] = 8'hF1;
DFS[16'h01AF] = 8'h20;
DFS[16'h01B0] = 8'h33;
DFS[16'h01B1] = 8'h80;
DFS[16'h01B2] = 8'hC8;
DFS[16'h01B3] = 8'h44;
DFS[16'h01B4] = 8'h69;
DFS[16'h01B5] = 8'h73;
DFS[16'h01B6] = 8'h6B;
DFS[16'h01B7] = 8'h20;
DFS[16'h01B8] = 8'h63;
DFS[16'h01B9] = 8'h68;
DFS[16'h01BA] = 8'h61;
DFS[16'h01BB] = 8'h6E;
DFS[16'h01BC] = 8'h67;
DFS[16'h01BD] = 8'h65;
DFS[16'h01BE] = 8'h64;
DFS[16'h01BF] = 8'h00;
DFS[16'h01C0] = 8'h20;
DFS[16'h01C1] = 8'hE1;
DFS[16'h01C2] = 8'h83;
DFS[16'h01C3] = 8'hB9;
DFS[16'h01C4] = 8'h0F;
DFS[16'h01C5] = 8'h0E;
DFS[16'h01C6] = 8'h08;
DFS[16'h01C7] = 8'h29;
DFS[16'h01C8] = 8'h7F;
DFS[16'h01C9] = 8'hD0;
DFS[16'h01CA] = 8'h05;
DFS[16'h01CB] = 8'h20;
DFS[16'h01CC] = 8'hCB;
DFS[16'h01CD] = 8'h9F;
DFS[16'h01CE] = 8'hF0;
DFS[16'h01CF] = 8'h06;
DFS[16'h01D0] = 8'h20;
DFS[16'h01D1] = 8'h9C;
DFS[16'h01D2] = 8'h80;
DFS[16'h01D3] = 8'h20;
DFS[16'h01D4] = 8'h9A;
DFS[16'h01D5] = 8'h80;
DFS[16'h01D6] = 8'hA2;
DFS[16'h01D7] = 8'h06;
DFS[16'h01D8] = 8'hB9;
DFS[16'h01D9] = 8'h08;
DFS[16'h01DA] = 8'h0E;
DFS[16'h01DB] = 8'h29;
DFS[16'h01DC] = 8'h7F;
DFS[16'h01DD] = 8'h20;
DFS[16'h01DE] = 8'h9C;
DFS[16'h01DF] = 8'h80;
DFS[16'h01E0] = 8'hC8;
DFS[16'h01E1] = 8'hCA;
DFS[16'h01E2] = 8'h10;
DFS[16'h01E3] = 8'hF4;
DFS[16'h01E4] = 8'h20;
DFS[16'h01E5] = 8'hCB;
DFS[16'h01E6] = 8'h9F;
DFS[16'h01E7] = 8'hA9;
DFS[16'h01E8] = 8'h20;
DFS[16'h01E9] = 8'h28;
DFS[16'h01EA] = 8'h10;
DFS[16'h01EB] = 8'h02;
DFS[16'h01EC] = 8'hA9;
DFS[16'h01ED] = 8'h4C;
DFS[16'h01EE] = 8'h20;
DFS[16'h01EF] = 8'h9C;
DFS[16'h01F0] = 8'h80;
DFS[16'h01F1] = 8'h4C;
DFS[16'h01F2] = 8'hCE;
DFS[16'h01F3] = 8'h9F;
DFS[16'h01F4] = 8'h20;
DFS[16'h01F5] = 8'hCE;
DFS[16'h01F6] = 8'h9F;
DFS[16'h01F7] = 8'h88;
DFS[16'h01F8] = 8'hD0;
DFS[16'h01F9] = 8'hFA;
DFS[16'h01FA] = 8'h60;
DFS[16'h01FB] = 8'h4A;
DFS[16'h01FC] = 8'h4A;
DFS[16'h01FD] = 8'h4A;
DFS[16'h01FE] = 8'h4A;
DFS[16'h01FF] = 8'h4A;
DFS[16'h0200] = 8'h4A;
DFS[16'h0201] = 8'h29;
DFS[16'h0202] = 8'h03;
DFS[16'h0203] = 8'h60;
DFS[16'h0204] = 8'h4A;
DFS[16'h0205] = 8'h4A;
DFS[16'h0206] = 8'h4A;
DFS[16'h0207] = 8'h4A;
DFS[16'h0208] = 8'h4A;
DFS[16'h0209] = 8'h60;
DFS[16'h020A] = 8'h0A;
DFS[16'h020B] = 8'h0A;
DFS[16'h020C] = 8'h0A;
DFS[16'h020D] = 8'h0A;
DFS[16'h020E] = 8'h0A;
DFS[16'h020F] = 8'h60;
DFS[16'h0210] = 8'hC8;
DFS[16'h0211] = 8'hC8;
DFS[16'h0212] = 8'hC8;
DFS[16'h0213] = 8'hC8;
DFS[16'h0214] = 8'hC8;
DFS[16'h0215] = 8'hC8;
DFS[16'h0216] = 8'hC8;
DFS[16'h0217] = 8'hC8;
DFS[16'h0218] = 8'h60;
DFS[16'h0219] = 8'h88;
DFS[16'h021A] = 8'h88;
DFS[16'h021B] = 8'h88;
DFS[16'h021C] = 8'h88;
DFS[16'h021D] = 8'h88;
DFS[16'h021E] = 8'h88;
DFS[16'h021F] = 8'h88;
DFS[16'h0220] = 8'h88;
DFS[16'h0221] = 8'h60;
DFS[16'h0222] = 8'h00;
DFS[16'h0223] = 8'h00;
DFS[16'h0224] = 8'h00;
DFS[16'h0225] = 8'h00;
DFS[16'h0226] = 8'h00;
DFS[16'h0227] = 8'h00;
DFS[16'h0228] = 8'h00;
DFS[16'h0229] = 8'h00;
DFS[16'h022A] = 8'h00;
DFS[16'h022B] = 8'h00;
DFS[16'h022C] = 8'h00;
DFS[16'h022D] = 8'h00;
DFS[16'h022E] = 8'h00;
DFS[16'h022F] = 8'h00;
DFS[16'h0230] = 8'h00;
DFS[16'h0231] = 8'h00;
DFS[16'h0232] = 8'h00;
DFS[16'h0233] = 8'h00;
DFS[16'h0234] = 8'h00;
DFS[16'h0235] = 8'h00;
DFS[16'h0236] = 8'h00;
DFS[16'h0237] = 8'h00;
DFS[16'h0238] = 8'h00;
DFS[16'h0239] = 8'h00;
DFS[16'h023A] = 8'h00;
DFS[16'h023B] = 8'h00;
DFS[16'h023C] = 8'h00;
DFS[16'h023D] = 8'h00;
DFS[16'h023E] = 8'h00;
DFS[16'h023F] = 8'h00;
DFS[16'h0240] = 8'h00;
DFS[16'h0241] = 8'h00;
DFS[16'h0242] = 8'h00;
DFS[16'h0243] = 8'h00;
DFS[16'h0244] = 8'h00;
DFS[16'h0245] = 8'h00;
DFS[16'h0246] = 8'h00;
DFS[16'h0247] = 8'h00;
DFS[16'h0248] = 8'h00;
DFS[16'h0249] = 8'h00;
DFS[16'h024A] = 8'h00;
DFS[16'h024B] = 8'h00;
DFS[16'h024C] = 8'h00;
DFS[16'h024D] = 8'h00;
DFS[16'h024E] = 8'h00;
DFS[16'h024F] = 8'h00;
DFS[16'h0250] = 8'h00;
DFS[16'h0251] = 8'h00;
DFS[16'h0252] = 8'h00;
DFS[16'h0253] = 8'h00;
DFS[16'h0254] = 8'h00;
DFS[16'h0255] = 8'h00;
DFS[16'h0256] = 8'h00;
DFS[16'h0257] = 8'h00;
DFS[16'h0258] = 8'h00;
DFS[16'h0259] = 8'h00;
DFS[16'h025A] = 8'h00;
DFS[16'h025B] = 8'h00;
DFS[16'h025C] = 8'h00;
DFS[16'h025D] = 8'h60;
DFS[16'h025E] = 8'hA9;
DFS[16'h025F] = 8'h23;
DFS[16'h0260] = 8'hD0;
DFS[16'h0261] = 8'h02;
DFS[16'h0262] = 8'hA9;
DFS[16'h0263] = 8'hFF;
DFS[16'h0264] = 8'h8D;
DFS[16'h0265] = 8'hCF;
DFS[16'h0266] = 8'h10;
DFS[16'h0267] = 8'h60;
DFS[16'h0268] = 8'h20;
DFS[16'h0269] = 8'hFE;
DFS[16'h026A] = 8'h80;
DFS[16'h026B] = 8'h4C;
DFS[16'h026C] = 8'h71;
DFS[16'h026D] = 8'h82;
DFS[16'h026E] = 8'h20;
DFS[16'h026F] = 8'h06;
DFS[16'h0270] = 8'h81;
DFS[16'h0271] = 8'h20;
DFS[16'h0272] = 8'h96;
DFS[16'h0273] = 8'h82;
DFS[16'h0274] = 8'hB0;
DFS[16'h0275] = 8'hE7;
DFS[16'h0276] = 8'h20;
DFS[16'h0277] = 8'h2B;
DFS[16'h0278] = 8'h80;
DFS[16'h0279] = 8'hD6;
DFS[16'h027A] = 8'h6E;
DFS[16'h027B] = 8'h6F;
DFS[16'h027C] = 8'h74;
DFS[16'h027D] = 8'h20;
DFS[16'h027E] = 8'h66;
DFS[16'h027F] = 8'h6F;
DFS[16'h0280] = 8'h75;
DFS[16'h0281] = 8'h6E;
DFS[16'h0282] = 8'h64;
DFS[16'h0283] = 8'h00;
DFS[16'h0284] = 8'h20;
DFS[16'h0285] = 8'h5E;
DFS[16'h0286] = 8'h82;
DFS[16'h0287] = 8'h20;
DFS[16'h0288] = 8'h01;
DFS[16'h0289] = 8'h9A;
DFS[16'h028A] = 8'h20;
DFS[16'h028B] = 8'h68;
DFS[16'h028C] = 8'h82;
DFS[16'h028D] = 8'h20;
DFS[16'h028E] = 8'h01;
DFS[16'h028F] = 8'h83;
DFS[16'h0290] = 8'h20;
DFS[16'h0291] = 8'h9D;
DFS[16'h0292] = 8'h82;
DFS[16'h0293] = 8'hB0;
DFS[16'h0294] = 8'hF8;
DFS[16'h0295] = 8'h60;
DFS[16'h0296] = 8'h20;
DFS[16'h0297] = 8'h4D;
DFS[16'h0298] = 8'hAB;
DFS[16'h0299] = 8'hA0;
DFS[16'h029A] = 8'hF8;
DFS[16'h029B] = 8'hD0;
DFS[16'h029C] = 8'h03;
DFS[16'h029D] = 8'hAC;
DFS[16'h029E] = 8'hCE;
DFS[16'h029F] = 8'h10;
DFS[16'h02A0] = 8'h20;
DFS[16'h02A1] = 8'h10;
DFS[16'h02A2] = 8'h82;
DFS[16'h02A3] = 8'hCC;
DFS[16'h02A4] = 8'h05;
DFS[16'h02A5] = 8'h0F;
DFS[16'h02A6] = 8'hB0;
DFS[16'h02A7] = 8'h44;
DFS[16'h02A8] = 8'h20;
DFS[16'h02A9] = 8'h10;
DFS[16'h02AA] = 8'h82;
DFS[16'h02AB] = 8'hA2;
DFS[16'h02AC] = 8'h07;
DFS[16'h02AD] = 8'hB5;
DFS[16'h02AE] = 8'hC7;
DFS[16'h02AF] = 8'hCD;
DFS[16'h02B0] = 8'hCF;
DFS[16'h02B1] = 8'h10;
DFS[16'h02B2] = 8'hF0;
DFS[16'h02B3] = 8'h0E;
DFS[16'h02B4] = 8'h20;
DFS[16'h02B5] = 8'hEE;
DFS[16'h02B6] = 8'h82;
DFS[16'h02B7] = 8'h59;
DFS[16'h02B8] = 8'h07;
DFS[16'h02B9] = 8'h0E;
DFS[16'h02BA] = 8'hB0;
DFS[16'h02BB] = 8'h02;
DFS[16'h02BC] = 8'h29;
DFS[16'h02BD] = 8'hDF;
DFS[16'h02BE] = 8'h29;
DFS[16'h02BF] = 8'h7F;
DFS[16'h02C0] = 8'hD0;
DFS[16'h02C1] = 8'h09;
DFS[16'h02C2] = 8'h88;
DFS[16'h02C3] = 8'hCA;
DFS[16'h02C4] = 8'h10;
DFS[16'h02C5] = 8'hE7;
DFS[16'h02C6] = 8'h8C;
DFS[16'h02C7] = 8'hCE;
DFS[16'h02C8] = 8'h10;
DFS[16'h02C9] = 8'h38;
DFS[16'h02CA] = 8'h60;
DFS[16'h02CB] = 8'h88;
DFS[16'h02CC] = 8'hCA;
DFS[16'h02CD] = 8'h10;
DFS[16'h02CE] = 8'hFC;
DFS[16'h02CF] = 8'h30;
DFS[16'h02D0] = 8'hCF;
DFS[16'h02D1] = 8'h20;
DFS[16'h02D2] = 8'h4C;
DFS[16'h02D3] = 8'h98;
DFS[16'h02D4] = 8'hB9;
DFS[16'h02D5] = 8'h10;
DFS[16'h02D6] = 8'h0E;
DFS[16'h02D7] = 8'h99;
DFS[16'h02D8] = 8'h08;
DFS[16'h02D9] = 8'h0E;
DFS[16'h02DA] = 8'hB9;
DFS[16'h02DB] = 8'h10;
DFS[16'h02DC] = 8'h0F;
DFS[16'h02DD] = 8'h99;
DFS[16'h02DE] = 8'h08;
DFS[16'h02DF] = 8'h0F;
DFS[16'h02E0] = 8'hC8;
DFS[16'h02E1] = 8'hCC;
DFS[16'h02E2] = 8'h05;
DFS[16'h02E3] = 8'h0F;
DFS[16'h02E4] = 8'h90;
DFS[16'h02E5] = 8'hEE;
DFS[16'h02E6] = 8'h98;
DFS[16'h02E7] = 8'hE9;
DFS[16'h02E8] = 8'h08;
DFS[16'h02E9] = 8'h8D;
DFS[16'h02EA] = 8'h05;
DFS[16'h02EB] = 8'h0F;
DFS[16'h02EC] = 8'h18;
DFS[16'h02ED] = 8'h60;
DFS[16'h02EE] = 8'h48;
DFS[16'h02EF] = 8'h29;
DFS[16'h02F0] = 8'hDF;
DFS[16'h02F1] = 8'hC9;
DFS[16'h02F2] = 8'h41;
DFS[16'h02F3] = 8'h90;
DFS[16'h02F4] = 8'h04;
DFS[16'h02F5] = 8'hC9;
DFS[16'h02F6] = 8'h5B;
DFS[16'h02F7] = 8'h90;
DFS[16'h02F8] = 8'h01;
DFS[16'h02F9] = 8'h38;
DFS[16'h02FA] = 8'h68;
DFS[16'h02FB] = 8'h60;
DFS[16'h02FC] = 8'h2C;
DFS[16'h02FD] = 8'hC7;
DFS[16'h02FE] = 8'h10;
DFS[16'h02FF] = 8'h30;
DFS[16'h0300] = 8'hEC;
DFS[16'h0301] = 8'h20;
DFS[16'h0302] = 8'hE1;
DFS[16'h0303] = 8'h83;
DFS[16'h0304] = 8'h20;
DFS[16'h0305] = 8'hC0;
DFS[16'h0306] = 8'h81;
DFS[16'h0307] = 8'h98;
DFS[16'h0308] = 8'h48;
DFS[16'h0309] = 8'hA9;
DFS[16'h030A] = 8'h60;
DFS[16'h030B] = 8'h85;
DFS[16'h030C] = 8'hB0;
DFS[16'h030D] = 8'hA9;
DFS[16'h030E] = 8'h10;
DFS[16'h030F] = 8'h85;
DFS[16'h0310] = 8'hB1;
DFS[16'h0311] = 8'h20;
DFS[16'h0312] = 8'h7E;
DFS[16'h0313] = 8'h83;
DFS[16'h0314] = 8'hA0;
DFS[16'h0315] = 8'h02;
DFS[16'h0316] = 8'h20;
DFS[16'h0317] = 8'hCE;
DFS[16'h0318] = 8'h9F;
DFS[16'h0319] = 8'h20;
DFS[16'h031A] = 8'h35;
DFS[16'h031B] = 8'h83;
DFS[16'h031C] = 8'h20;
DFS[16'h031D] = 8'h35;
DFS[16'h031E] = 8'h83;
DFS[16'h031F] = 8'h20;
DFS[16'h0320] = 8'h35;
DFS[16'h0321] = 8'h83;
DFS[16'h0322] = 8'h68;
DFS[16'h0323] = 8'hA8;
DFS[16'h0324] = 8'hB9;
DFS[16'h0325] = 8'h0E;
DFS[16'h0326] = 8'h0F;
DFS[16'h0327] = 8'h29;
DFS[16'h0328] = 8'h03;
DFS[16'h0329] = 8'h20;
DFS[16'h032A] = 8'hCA;
DFS[16'h032B] = 8'h80;
DFS[16'h032C] = 8'hB9;
DFS[16'h032D] = 8'h0F;
DFS[16'h032E] = 8'h0F;
DFS[16'h032F] = 8'h20;
DFS[16'h0330] = 8'hC2;
DFS[16'h0331] = 8'h80;
DFS[16'h0332] = 8'h4C;
DFS[16'h0333] = 8'h9A;
DFS[16'h0334] = 8'h9F;
DFS[16'h0335] = 8'hA2;
DFS[16'h0336] = 8'h03;
DFS[16'h0337] = 8'hB9;
DFS[16'h0338] = 8'h62;
DFS[16'h0339] = 8'h10;
DFS[16'h033A] = 8'h20;
DFS[16'h033B] = 8'hC2;
DFS[16'h033C] = 8'h80;
DFS[16'h033D] = 8'h88;
DFS[16'h033E] = 8'hCA;
DFS[16'h033F] = 8'hD0;
DFS[16'h0340] = 8'hF6;
DFS[16'h0341] = 8'h20;
DFS[16'h0342] = 8'h11;
DFS[16'h0343] = 8'h82;
DFS[16'h0344] = 8'h4C;
DFS[16'h0345] = 8'hCE;
DFS[16'h0346] = 8'h9F;
DFS[16'h0347] = 8'h20;
DFS[16'h0348] = 8'hE1;
DFS[16'h0349] = 8'h83;
DFS[16'h034A] = 8'h4C;
DFS[16'h034B] = 8'h4D;
DFS[16'h034C] = 8'hAB;
DFS[16'h034D] = 8'hAD;
DFS[16'h034E] = 8'hCA;
DFS[16'h034F] = 8'h10;
DFS[16'h0350] = 8'h85;
DFS[16'h0351] = 8'hCE;
DFS[16'h0352] = 8'hAD;
DFS[16'h0353] = 8'hCB;
DFS[16'h0354] = 8'h10;
DFS[16'h0355] = 8'h4C;
DFS[16'h0356] = 8'h7E;
DFS[16'h0357] = 8'h87;
DFS[16'h0358] = 8'h20;
DFS[16'h0359] = 8'hBF;
DFS[16'h035A] = 8'h86;
DFS[16'h035B] = 8'hF0;
DFS[16'h035C] = 8'hF5;
DFS[16'h035D] = 8'h20;
DFS[16'h035E] = 8'hC5;
DFS[16'h035F] = 8'hFF;
DFS[16'h0360] = 8'hB0;
DFS[16'h0361] = 8'h12;
DFS[16'h0362] = 8'hC9;
DFS[16'h0363] = 8'h3A;
DFS[16'h0364] = 8'hF0;
DFS[16'h0365] = 8'hF7;
DFS[16'h0366] = 8'h38;
DFS[16'h0367] = 8'hE9;
DFS[16'h0368] = 8'h30;
DFS[16'h0369] = 8'h90;
DFS[16'h036A] = 8'h09;
DFS[16'h036B] = 8'hC9;
DFS[16'h036C] = 8'h04;
DFS[16'h036D] = 8'hB0;
DFS[16'h036E] = 8'h05;
DFS[16'h036F] = 8'h20;
DFS[16'h0370] = 8'h7E;
DFS[16'h0371] = 8'h87;
DFS[16'h0372] = 8'h18;
DFS[16'h0373] = 8'h60;
DFS[16'h0374] = 8'h20;
DFS[16'h0375] = 8'h22;
DFS[16'h0376] = 8'h80;
DFS[16'h0377] = 8'hCD;
DFS[16'h0378] = 8'h64;
DFS[16'h0379] = 8'h72;
DFS[16'h037A] = 8'h69;
DFS[16'h037B] = 8'h76;
DFS[16'h037C] = 8'h65;
DFS[16'h037D] = 8'h00;
DFS[16'h037E] = 8'h20;
DFS[16'h037F] = 8'hE1;
DFS[16'h0380] = 8'h83;
DFS[16'h0381] = 8'h98;
DFS[16'h0382] = 8'h48;
DFS[16'h0383] = 8'hAA;
DFS[16'h0384] = 8'hA0;
DFS[16'h0385] = 8'h02;
DFS[16'h0386] = 8'hA9;
DFS[16'h0387] = 8'h00;
DFS[16'h0388] = 8'h91;
DFS[16'h0389] = 8'hB0;
DFS[16'h038A] = 8'hC8;
DFS[16'h038B] = 8'hC0;
DFS[16'h038C] = 8'h12;
DFS[16'h038D] = 8'hD0;
DFS[16'h038E] = 8'hF9;
DFS[16'h038F] = 8'hA0;
DFS[16'h0390] = 8'h02;
DFS[16'h0391] = 8'h20;
DFS[16'h0392] = 8'hCF;
DFS[16'h0393] = 8'h83;
DFS[16'h0394] = 8'hC8;
DFS[16'h0395] = 8'hC8;
DFS[16'h0396] = 8'hC0;
DFS[16'h0397] = 8'h0E;
DFS[16'h0398] = 8'hD0;
DFS[16'h0399] = 8'hF7;
DFS[16'h039A] = 8'h68;
DFS[16'h039B] = 8'hAA;
DFS[16'h039C] = 8'hBD;
DFS[16'h039D] = 8'h0F;
DFS[16'h039E] = 8'h0E;
DFS[16'h039F] = 8'h10;
DFS[16'h03A0] = 8'h06;
DFS[16'h03A1] = 8'hA9;
DFS[16'h03A2] = 8'h0A;
DFS[16'h03A3] = 8'hA0;
DFS[16'h03A4] = 8'h0E;
DFS[16'h03A5] = 8'h91;
DFS[16'h03A6] = 8'hB0;
DFS[16'h03A7] = 8'hBD;
DFS[16'h03A8] = 8'h0E;
DFS[16'h03A9] = 8'h0F;
DFS[16'h03AA] = 8'hA0;
DFS[16'h03AB] = 8'h04;
DFS[16'h03AC] = 8'h20;
DFS[16'h03AD] = 8'hBB;
DFS[16'h03AE] = 8'h83;
DFS[16'h03AF] = 8'hA0;
DFS[16'h03B0] = 8'h0C;
DFS[16'h03B1] = 8'h4A;
DFS[16'h03B2] = 8'h4A;
DFS[16'h03B3] = 8'h48;
DFS[16'h03B4] = 8'h29;
DFS[16'h03B5] = 8'h03;
DFS[16'h03B6] = 8'h91;
DFS[16'h03B7] = 8'hB0;
DFS[16'h03B8] = 8'h68;
DFS[16'h03B9] = 8'hA0;
DFS[16'h03BA] = 8'h08;
DFS[16'h03BB] = 8'h4A;
DFS[16'h03BC] = 8'h4A;
DFS[16'h03BD] = 8'h48;
DFS[16'h03BE] = 8'h29;
DFS[16'h03BF] = 8'h03;
DFS[16'h03C0] = 8'h91;
DFS[16'h03C1] = 8'hB0;
DFS[16'h03C2] = 8'hC9;
DFS[16'h03C3] = 8'h03;
DFS[16'h03C4] = 8'hD0;
DFS[16'h03C5] = 8'h07;
DFS[16'h03C6] = 8'hA9;
DFS[16'h03C7] = 8'hFF;
DFS[16'h03C8] = 8'h91;
DFS[16'h03C9] = 8'hB0;
DFS[16'h03CA] = 8'hC8;
DFS[16'h03CB] = 8'h91;
DFS[16'h03CC] = 8'hB0;
DFS[16'h03CD] = 8'h68;
DFS[16'h03CE] = 8'h60;
DFS[16'h03CF] = 8'h20;
DFS[16'h03D0] = 8'hD2;
DFS[16'h03D1] = 8'h83;
DFS[16'h03D2] = 8'hBD;
DFS[16'h03D3] = 8'h08;
DFS[16'h03D4] = 8'h0F;
DFS[16'h03D5] = 8'h91;
DFS[16'h03D6] = 8'hB0;
DFS[16'h03D7] = 8'hE8;
DFS[16'h03D8] = 8'hC8;
DFS[16'h03D9] = 8'h60;
DFS[16'h03DA] = 8'hE6;
DFS[16'h03DB] = 8'hAE;
DFS[16'h03DC] = 8'hD0;
DFS[16'h03DD] = 8'h02;
DFS[16'h03DE] = 8'hE6;
DFS[16'h03DF] = 8'hAF;
DFS[16'h03E0] = 8'h60;
DFS[16'h03E1] = 8'h48;
DFS[16'h03E2] = 8'h8A;
DFS[16'h03E3] = 8'h48;
DFS[16'h03E4] = 8'h98;
DFS[16'h03E5] = 8'h48;
DFS[16'h03E6] = 8'hA9;
DFS[16'h03E7] = 8'h84;
DFS[16'h03E8] = 8'h48;
DFS[16'h03E9] = 8'hA9;
DFS[16'h03EA] = 8'h03;
DFS[16'h03EB] = 8'h48;
DFS[16'h03EC] = 8'hA0;
DFS[16'h03ED] = 8'h05;
DFS[16'h03EE] = 8'hBA;
DFS[16'h03EF] = 8'hBD;
DFS[16'h03F0] = 8'h07;
DFS[16'h03F1] = 8'h01;
DFS[16'h03F2] = 8'h48;
DFS[16'h03F3] = 8'h88;
DFS[16'h03F4] = 8'hD0;
DFS[16'h03F5] = 8'hF8;
DFS[16'h03F6] = 8'hA0;
DFS[16'h03F7] = 8'h0A;
DFS[16'h03F8] = 8'hBD;
DFS[16'h03F9] = 8'h09;
DFS[16'h03FA] = 8'h01;
DFS[16'h03FB] = 8'h9D;
DFS[16'h03FC] = 8'h0B;
DFS[16'h03FD] = 8'h01;
DFS[16'h03FE] = 8'hCA;
DFS[16'h03FF] = 8'h88;
DFS[16'h0400] = 8'hD0;
DFS[16'h0401] = 8'hF6;
DFS[16'h0402] = 8'h68;
DFS[16'h0403] = 8'h68;
DFS[16'h0404] = 8'h68;
DFS[16'h0405] = 8'hA8;
DFS[16'h0406] = 8'h68;
DFS[16'h0407] = 8'hAA;
DFS[16'h0408] = 8'h68;
DFS[16'h0409] = 8'h60;
DFS[16'h040A] = 8'hBA;
DFS[16'h040B] = 8'h9D;
DFS[16'h040C] = 8'h03;
DFS[16'h040D] = 8'h01;
DFS[16'h040E] = 8'h4C;
DFS[16'h040F] = 8'h04;
DFS[16'h0410] = 8'h84;
DFS[16'h0411] = 8'h48;
DFS[16'h0412] = 8'h8A;
DFS[16'h0413] = 8'h48;
DFS[16'h0414] = 8'h98;
DFS[16'h0415] = 8'h48;
DFS[16'h0416] = 8'hA9;
DFS[16'h0417] = 8'h84;
DFS[16'h0418] = 8'h48;
DFS[16'h0419] = 8'hA9;
DFS[16'h041A] = 8'h09;
DFS[16'h041B] = 8'h48;
DFS[16'h041C] = 8'hD0;
DFS[16'h041D] = 8'hCE;
DFS[16'h041E] = 8'h20;
DFS[16'h041F] = 8'hB8;
DFS[16'h0420] = 8'h86;
DFS[16'h0421] = 8'h20;
DFS[16'h0422] = 8'h47;
DFS[16'h0423] = 8'hAB;
DFS[16'h0424] = 8'hA0;
DFS[16'h0425] = 8'hFF;
DFS[16'h0426] = 8'h84;
DFS[16'h0427] = 8'hA8;
DFS[16'h0428] = 8'hC8;
DFS[16'h0429] = 8'h84;
DFS[16'h042A] = 8'hAA;
DFS[16'h042B] = 8'hB9;
DFS[16'h042C] = 8'h00;
DFS[16'h042D] = 8'h0E;
DFS[16'h042E] = 8'hC0;
DFS[16'h042F] = 8'h08;
DFS[16'h0430] = 8'h90;
DFS[16'h0431] = 8'h03;
DFS[16'h0432] = 8'hB9;
DFS[16'h0433] = 8'hF8;
DFS[16'h0434] = 8'h0E;
DFS[16'h0435] = 8'h20;
DFS[16'h0436] = 8'h9C;
DFS[16'h0437] = 8'h80;
DFS[16'h0438] = 8'hC8;
DFS[16'h0439] = 8'hC0;
DFS[16'h043A] = 8'h0C;
DFS[16'h043B] = 8'hD0;
DFS[16'h043C] = 8'hEE;
DFS[16'h043D] = 8'h20;
DFS[16'h043E] = 8'h65;
DFS[16'h043F] = 8'h80;
DFS[16'h0440] = 8'h20;
DFS[16'h0441] = 8'h28;
DFS[16'h0442] = 8'hAD;
DFS[16'h0443] = 8'h04;
DFS[16'h0444] = 8'h0F;
DFS[16'h0445] = 8'h20;
DFS[16'h0446] = 8'hC2;
DFS[16'h0447] = 8'h80;
DFS[16'h0448] = 8'h20;
DFS[16'h0449] = 8'h65;
DFS[16'h044A] = 8'h80;
DFS[16'h044B] = 8'h29;
DFS[16'h044C] = 8'h0D;
DFS[16'h044D] = 8'h44;
DFS[16'h044E] = 8'h72;
DFS[16'h044F] = 8'h69;
DFS[16'h0450] = 8'h76;
DFS[16'h0451] = 8'h65;
DFS[16'h0452] = 8'h20;
DFS[16'h0453] = 8'hA5;
DFS[16'h0454] = 8'hCF;
DFS[16'h0455] = 8'h20;
DFS[16'h0456] = 8'hCA;
DFS[16'h0457] = 8'h80;
DFS[16'h0458] = 8'hA0;
DFS[16'h0459] = 8'h0D;
DFS[16'h045A] = 8'h20;
DFS[16'h045B] = 8'hF4;
DFS[16'h045C] = 8'h81;
DFS[16'h045D] = 8'h20;
DFS[16'h045E] = 8'h65;
DFS[16'h045F] = 8'h80;
DFS[16'h0460] = 8'h4F;
DFS[16'h0461] = 8'h70;
DFS[16'h0462] = 8'h74;
DFS[16'h0463] = 8'h69;
DFS[16'h0464] = 8'h6F;
DFS[16'h0465] = 8'h6E;
DFS[16'h0466] = 8'h20;
DFS[16'h0467] = 8'hAD;
DFS[16'h0468] = 8'h06;
DFS[16'h0469] = 8'h0F;
DFS[16'h046A] = 8'h20;
DFS[16'h046B] = 8'h05;
DFS[16'h046C] = 8'h82;
DFS[16'h046D] = 8'h20;
DFS[16'h046E] = 8'hCA;
DFS[16'h046F] = 8'h80;
DFS[16'h0470] = 8'h20;
DFS[16'h0471] = 8'h65;
DFS[16'h0472] = 8'h80;
DFS[16'h0473] = 8'h20;
DFS[16'h0474] = 8'h28;
DFS[16'h0475] = 8'hA0;
DFS[16'h0476] = 8'h03;
DFS[16'h0477] = 8'h0A;
DFS[16'h0478] = 8'h0A;
DFS[16'h0479] = 8'hAA;
DFS[16'h047A] = 8'hBD;
DFS[16'h047B] = 8'h6F;
DFS[16'h047C] = 8'h85;
DFS[16'h047D] = 8'h20;
DFS[16'h047E] = 8'h9C;
DFS[16'h047F] = 8'h80;
DFS[16'h0480] = 8'hE8;
DFS[16'h0481] = 8'h88;
DFS[16'h0482] = 8'h10;
DFS[16'h0483] = 8'hF6;
DFS[16'h0484] = 8'h20;
DFS[16'h0485] = 8'h65;
DFS[16'h0486] = 8'h80;
DFS[16'h0487] = 8'h29;
DFS[16'h0488] = 8'h0D;
DFS[16'h0489] = 8'h44;
DFS[16'h048A] = 8'h69;
DFS[16'h048B] = 8'h72;
DFS[16'h048C] = 8'h65;
DFS[16'h048D] = 8'h63;
DFS[16'h048E] = 8'h74;
DFS[16'h048F] = 8'h6F;
DFS[16'h0490] = 8'h72;
DFS[16'h0491] = 8'h79;
DFS[16'h0492] = 8'h20;
DFS[16'h0493] = 8'h3A;
DFS[16'h0494] = 8'hAD;
DFS[16'h0495] = 8'hCB;
DFS[16'h0496] = 8'h10;
DFS[16'h0497] = 8'h20;
DFS[16'h0498] = 8'hCA;
DFS[16'h0499] = 8'h80;
DFS[16'h049A] = 8'h20;
DFS[16'h049B] = 8'h9A;
DFS[16'h049C] = 8'h80;
DFS[16'h049D] = 8'hAD;
DFS[16'h049E] = 8'hCA;
DFS[16'h049F] = 8'h10;
DFS[16'h04A0] = 8'h20;
DFS[16'h04A1] = 8'h9C;
DFS[16'h04A2] = 8'h80;
DFS[16'h04A3] = 8'hA0;
DFS[16'h04A4] = 8'h06;
DFS[16'h04A5] = 8'h20;
DFS[16'h04A6] = 8'hF4;
DFS[16'h04A7] = 8'h81;
DFS[16'h04A8] = 8'h20;
DFS[16'h04A9] = 8'h65;
DFS[16'h04AA] = 8'h80;
DFS[16'h04AB] = 8'h4C;
DFS[16'h04AC] = 8'h69;
DFS[16'h04AD] = 8'h62;
DFS[16'h04AE] = 8'h72;
DFS[16'h04AF] = 8'h61;
DFS[16'h04B0] = 8'h72;
DFS[16'h04B1] = 8'h79;
DFS[16'h04B2] = 8'h20;
DFS[16'h04B3] = 8'h3A;
DFS[16'h04B4] = 8'hAD;
DFS[16'h04B5] = 8'hCD;
DFS[16'h04B6] = 8'h10;
DFS[16'h04B7] = 8'h20;
DFS[16'h04B8] = 8'hCA;
DFS[16'h04B9] = 8'h80;
DFS[16'h04BA] = 8'h20;
DFS[16'h04BB] = 8'h9A;
DFS[16'h04BC] = 8'h80;
DFS[16'h04BD] = 8'hAD;
DFS[16'h04BE] = 8'hCC;
DFS[16'h04BF] = 8'h10;
DFS[16'h04C0] = 8'h20;
DFS[16'h04C1] = 8'h9C;
DFS[16'h04C2] = 8'h80;
DFS[16'h04C3] = 8'h20;
DFS[16'h04C4] = 8'h9A;
DFS[16'h04C5] = 8'h9F;
DFS[16'h04C6] = 8'hA0;
DFS[16'h04C7] = 8'h00;
DFS[16'h04C8] = 8'hCC;
DFS[16'h04C9] = 8'h05;
DFS[16'h04CA] = 8'h0F;
DFS[16'h04CB] = 8'hB0;
DFS[16'h04CC] = 8'h17;
DFS[16'h04CD] = 8'hB9;
DFS[16'h04CE] = 8'h0F;
DFS[16'h04CF] = 8'h0E;
DFS[16'h04D0] = 8'h4D;
DFS[16'h04D1] = 8'hCA;
DFS[16'h04D2] = 8'h10;
DFS[16'h04D3] = 8'h29;
DFS[16'h04D4] = 8'h7F;
DFS[16'h04D5] = 8'hD0;
DFS[16'h04D6] = 8'h08;
DFS[16'h04D7] = 8'hB9;
DFS[16'h04D8] = 8'h0F;
DFS[16'h04D9] = 8'h0E;
DFS[16'h04DA] = 8'h29;
DFS[16'h04DB] = 8'h80;
DFS[16'h04DC] = 8'h99;
DFS[16'h04DD] = 8'h0F;
DFS[16'h04DE] = 8'h0E;
DFS[16'h04DF] = 8'h20;
DFS[16'h04E0] = 8'h10;
DFS[16'h04E1] = 8'h82;
DFS[16'h04E2] = 8'h90;
DFS[16'h04E3] = 8'hE4;
DFS[16'h04E4] = 8'hA0;
DFS[16'h04E5] = 8'h00;
DFS[16'h04E6] = 8'h20;
DFS[16'h04E7] = 8'hF6;
DFS[16'h04E8] = 8'h84;
DFS[16'h04E9] = 8'h90;
DFS[16'h04EA] = 8'h16;
DFS[16'h04EB] = 8'hA9;
DFS[16'h04EC] = 8'hFF;
DFS[16'h04ED] = 8'h8D;
DFS[16'h04EE] = 8'h82;
DFS[16'h04EF] = 8'h10;
DFS[16'h04F0] = 8'h4C;
DFS[16'h04F1] = 8'h9A;
DFS[16'h04F2] = 8'h9F;
DFS[16'h04F3] = 8'h20;
DFS[16'h04F4] = 8'h10;
DFS[16'h04F5] = 8'h82;
DFS[16'h04F6] = 8'hCC;
DFS[16'h04F7] = 8'h05;
DFS[16'h04F8] = 8'h0F;
DFS[16'h04F9] = 8'hB0;
DFS[16'h04FA] = 8'h05;
DFS[16'h04FB] = 8'hB9;
DFS[16'h04FC] = 8'h08;
DFS[16'h04FD] = 8'h0E;
DFS[16'h04FE] = 8'h30;
DFS[16'h04FF] = 8'hF3;
DFS[16'h0500] = 8'h60;
DFS[16'h0501] = 8'h84;
DFS[16'h0502] = 8'hAB;
DFS[16'h0503] = 8'hA2;
DFS[16'h0504] = 8'h00;
DFS[16'h0505] = 8'hB9;
DFS[16'h0506] = 8'h08;
DFS[16'h0507] = 8'h0E;
DFS[16'h0508] = 8'h29;
DFS[16'h0509] = 8'h7F;
DFS[16'h050A] = 8'h9D;
DFS[16'h050B] = 8'h60;
DFS[16'h050C] = 8'h10;
DFS[16'h050D] = 8'hC8;
DFS[16'h050E] = 8'hE8;
DFS[16'h050F] = 8'hE0;
DFS[16'h0510] = 8'h08;
DFS[16'h0511] = 8'hD0;
DFS[16'h0512] = 8'hF2;
DFS[16'h0513] = 8'h20;
DFS[16'h0514] = 8'hF6;
DFS[16'h0515] = 8'h84;
DFS[16'h0516] = 8'hB0;
DFS[16'h0517] = 8'h1F;
DFS[16'h0518] = 8'h38;
DFS[16'h0519] = 8'hA2;
DFS[16'h051A] = 8'h06;
DFS[16'h051B] = 8'hB9;
DFS[16'h051C] = 8'h0E;
DFS[16'h051D] = 8'h0E;
DFS[16'h051E] = 8'hFD;
DFS[16'h051F] = 8'h60;
DFS[16'h0520] = 8'h10;
DFS[16'h0521] = 8'h88;
DFS[16'h0522] = 8'hCA;
DFS[16'h0523] = 8'h10;
DFS[16'h0524] = 8'hF6;
DFS[16'h0525] = 8'h20;
DFS[16'h0526] = 8'h11;
DFS[16'h0527] = 8'h82;
DFS[16'h0528] = 8'hB9;
DFS[16'h0529] = 8'h0F;
DFS[16'h052A] = 8'h0E;
DFS[16'h052B] = 8'h29;
DFS[16'h052C] = 8'h7F;
DFS[16'h052D] = 8'hED;
DFS[16'h052E] = 8'h67;
DFS[16'h052F] = 8'h10;
DFS[16'h0530] = 8'h90;
DFS[16'h0531] = 8'hCF;
DFS[16'h0532] = 8'h20;
DFS[16'h0533] = 8'h10;
DFS[16'h0534] = 8'h82;
DFS[16'h0535] = 8'hB0;
DFS[16'h0536] = 8'hDC;
DFS[16'h0537] = 8'hA4;
DFS[16'h0538] = 8'hAB;
DFS[16'h0539] = 8'hB9;
DFS[16'h053A] = 8'h08;
DFS[16'h053B] = 8'h0E;
DFS[16'h053C] = 8'h09;
DFS[16'h053D] = 8'h80;
DFS[16'h053E] = 8'h99;
DFS[16'h053F] = 8'h08;
DFS[16'h0540] = 8'h0E;
DFS[16'h0541] = 8'hAD;
DFS[16'h0542] = 8'h67;
DFS[16'h0543] = 8'h10;
DFS[16'h0544] = 8'hC5;
DFS[16'h0545] = 8'hAA;
DFS[16'h0546] = 8'hF0;
DFS[16'h0547] = 8'h10;
DFS[16'h0548] = 8'hA6;
DFS[16'h0549] = 8'hAA;
DFS[16'h054A] = 8'h85;
DFS[16'h054B] = 8'hAA;
DFS[16'h054C] = 8'hD0;
DFS[16'h054D] = 8'h0A;
DFS[16'h054E] = 8'h20;
DFS[16'h054F] = 8'h9A;
DFS[16'h0550] = 8'h9F;
DFS[16'h0551] = 8'h20;
DFS[16'h0552] = 8'h9A;
DFS[16'h0553] = 8'h9F;
DFS[16'h0554] = 8'hA0;
DFS[16'h0555] = 8'hFF;
DFS[16'h0556] = 8'hD0;
DFS[16'h0557] = 8'h09;
DFS[16'h0558] = 8'hA4;
DFS[16'h0559] = 8'hA8;
DFS[16'h055A] = 8'hD0;
DFS[16'h055B] = 8'hF5;
DFS[16'h055C] = 8'hA0;
DFS[16'h055D] = 8'h05;
DFS[16'h055E] = 8'h20;
DFS[16'h055F] = 8'hF4;
DFS[16'h0560] = 8'h81;
DFS[16'h0561] = 8'hC8;
DFS[16'h0562] = 8'h84;
DFS[16'h0563] = 8'hA8;
DFS[16'h0564] = 8'hA4;
DFS[16'h0565] = 8'hAB;
DFS[16'h0566] = 8'h20;
DFS[16'h0567] = 8'hCB;
DFS[16'h0568] = 8'h9F;
DFS[16'h0569] = 8'h20;
DFS[16'h056A] = 8'hC0;
DFS[16'h056B] = 8'h81;
DFS[16'h056C] = 8'h4C;
DFS[16'h056D] = 8'hE4;
DFS[16'h056E] = 8'h84;
DFS[16'h056F] = 8'h6F;
DFS[16'h0570] = 8'h66;
DFS[16'h0571] = 8'h66;
DFS[16'h0572] = 8'h00;
DFS[16'h0573] = 8'h4C;
DFS[16'h0574] = 8'h4F;
DFS[16'h0575] = 8'h41;
DFS[16'h0576] = 8'h44;
DFS[16'h0577] = 8'h52;
DFS[16'h0578] = 8'h55;
DFS[16'h0579] = 8'h4E;
DFS[16'h057A] = 8'h00;
DFS[16'h057B] = 8'h45;
DFS[16'h057C] = 8'h58;
DFS[16'h057D] = 8'h45;
DFS[16'h057E] = 8'h43;
DFS[16'h057F] = 8'hB9;
DFS[16'h0580] = 8'h0E;
DFS[16'h0581] = 8'h0F;
DFS[16'h0582] = 8'h20;
DFS[16'h0583] = 8'hFD;
DFS[16'h0584] = 8'h81;
DFS[16'h0585] = 8'h85;
DFS[16'h0586] = 8'hC4;
DFS[16'h0587] = 8'h18;
DFS[16'h0588] = 8'hA9;
DFS[16'h0589] = 8'hFF;
DFS[16'h058A] = 8'h79;
DFS[16'h058B] = 8'h0C;
DFS[16'h058C] = 8'h0F;
DFS[16'h058D] = 8'hB9;
DFS[16'h058E] = 8'h0F;
DFS[16'h058F] = 8'h0F;
DFS[16'h0590] = 8'h79;
DFS[16'h0591] = 8'h0D;
DFS[16'h0592] = 8'h0F;
DFS[16'h0593] = 8'h85;
DFS[16'h0594] = 8'hC5;
DFS[16'h0595] = 8'hB9;
DFS[16'h0596] = 8'h0E;
DFS[16'h0597] = 8'h0F;
DFS[16'h0598] = 8'h29;
DFS[16'h0599] = 8'h03;
DFS[16'h059A] = 8'h65;
DFS[16'h059B] = 8'hC4;
DFS[16'h059C] = 8'h85;
DFS[16'h059D] = 8'hC4;
DFS[16'h059E] = 8'h38;
DFS[16'h059F] = 8'hB9;
DFS[16'h05A0] = 8'h07;
DFS[16'h05A1] = 8'h0F;
DFS[16'h05A2] = 8'hE5;
DFS[16'h05A3] = 8'hC5;
DFS[16'h05A4] = 8'h48;
DFS[16'h05A5] = 8'hB9;
DFS[16'h05A6] = 8'h06;
DFS[16'h05A7] = 8'h0F;
DFS[16'h05A8] = 8'h29;
DFS[16'h05A9] = 8'h03;
DFS[16'h05AA] = 8'hE5;
DFS[16'h05AB] = 8'hC4;
DFS[16'h05AC] = 8'hAA;
DFS[16'h05AD] = 8'hA9;
DFS[16'h05AE] = 8'h00;
DFS[16'h05AF] = 8'hC5;
DFS[16'h05B0] = 8'hC2;
DFS[16'h05B1] = 8'h68;
DFS[16'h05B2] = 8'hE5;
DFS[16'h05B3] = 8'hC3;
DFS[16'h05B4] = 8'h8A;
DFS[16'h05B5] = 8'hE5;
DFS[16'h05B6] = 8'hC6;
DFS[16'h05B7] = 8'h60;
DFS[16'h05B8] = 8'h41;
DFS[16'h05B9] = 8'h43;
DFS[16'h05BA] = 8'h43;
DFS[16'h05BB] = 8'h45;
DFS[16'h05BC] = 8'h53;
DFS[16'h05BD] = 8'h53;
DFS[16'h05BE] = 8'h88;
DFS[16'h05BF] = 8'hD1;
DFS[16'h05C0] = 8'h32;
DFS[16'h05C1] = 8'h42;
DFS[16'h05C2] = 8'h41;
DFS[16'h05C3] = 8'h43;
DFS[16'h05C4] = 8'h4B;
DFS[16'h05C5] = 8'h55;
DFS[16'h05C6] = 8'h50;
DFS[16'h05C7] = 8'h9C;
DFS[16'h05C8] = 8'hBA;
DFS[16'h05C9] = 8'h54;
DFS[16'h05CA] = 8'h43;
DFS[16'h05CB] = 8'h4F;
DFS[16'h05CC] = 8'h4D;
DFS[16'h05CD] = 8'h50;
DFS[16'h05CE] = 8'h41;
DFS[16'h05CF] = 8'h43;
DFS[16'h05D0] = 8'h54;
DFS[16'h05D1] = 8'h9A;
DFS[16'h05D2] = 8'hBF;
DFS[16'h05D3] = 8'h0A;
DFS[16'h05D4] = 8'h43;
DFS[16'h05D5] = 8'h4F;
DFS[16'h05D6] = 8'h50;
DFS[16'h05D7] = 8'h59;
DFS[16'h05D8] = 8'h9D;
DFS[16'h05D9] = 8'h26;
DFS[16'h05DA] = 8'h64;
DFS[16'h05DB] = 8'h44;
DFS[16'h05DC] = 8'h45;
DFS[16'h05DD] = 8'h4C;
DFS[16'h05DE] = 8'h45;
DFS[16'h05DF] = 8'h54;
DFS[16'h05E0] = 8'h45;
DFS[16'h05E1] = 8'h86;
DFS[16'h05E2] = 8'hFD;
DFS[16'h05E3] = 8'h01;
DFS[16'h05E4] = 8'h44;
DFS[16'h05E5] = 8'h45;
DFS[16'h05E6] = 8'h53;
DFS[16'h05E7] = 8'h54;
DFS[16'h05E8] = 8'h52;
DFS[16'h05E9] = 8'h4F;
DFS[16'h05EA] = 8'h59;
DFS[16'h05EB] = 8'h87;
DFS[16'h05EC] = 8'h0F;
DFS[16'h05ED] = 8'h02;
DFS[16'h05EE] = 8'h44;
DFS[16'h05EF] = 8'h49;
DFS[16'h05F0] = 8'h52;
DFS[16'h05F1] = 8'h88;
DFS[16'h05F2] = 8'h4D;
DFS[16'h05F3] = 8'h09;
DFS[16'h05F4] = 8'h44;
DFS[16'h05F5] = 8'h52;
DFS[16'h05F6] = 8'h49;
DFS[16'h05F7] = 8'h56;
DFS[16'h05F8] = 8'h45;
DFS[16'h05F9] = 8'h87;
DFS[16'h05FA] = 8'h74;
DFS[16'h05FB] = 8'h0A;
DFS[16'h05FC] = 8'h45;
DFS[16'h05FD] = 8'h4E;
DFS[16'h05FE] = 8'h41;
DFS[16'h05FF] = 8'h42;
DFS[16'h0600] = 8'h4C;
DFS[16'h0601] = 8'h45;
DFS[16'h0602] = 8'h8A;
DFS[16'h0603] = 8'h38;
DFS[16'h0604] = 8'h00;
DFS[16'h0605] = 8'h49;
DFS[16'h0606] = 8'h4E;
DFS[16'h0607] = 8'h46;
DFS[16'h0608] = 8'h4F;
DFS[16'h0609] = 8'h82;
DFS[16'h060A] = 8'h83;
DFS[16'h060B] = 8'h02;
DFS[16'h060C] = 8'h4C;
DFS[16'h060D] = 8'h49;
DFS[16'h060E] = 8'h42;
DFS[16'h060F] = 8'h88;
DFS[16'h0610] = 8'h51;
DFS[16'h0611] = 8'h09;
DFS[16'h0612] = 8'h52;
DFS[16'h0613] = 8'h45;
DFS[16'h0614] = 8'h4E;
DFS[16'h0615] = 8'h41;
DFS[16'h0616] = 8'h4D;
DFS[16'h0617] = 8'h45;
DFS[16'h0618] = 8'h8A;
DFS[16'h0619] = 8'h6C;
DFS[16'h061A] = 8'h87;
DFS[16'h061B] = 8'h54;
DFS[16'h061C] = 8'h49;
DFS[16'h061D] = 8'h54;
DFS[16'h061E] = 8'h4C;
DFS[16'h061F] = 8'h45;
DFS[16'h0620] = 8'h88;
DFS[16'h0621] = 8'hA2;
DFS[16'h0622] = 8'h0B;
DFS[16'h0623] = 8'h57;
DFS[16'h0624] = 8'h49;
DFS[16'h0625] = 8'h50;
DFS[16'h0626] = 8'h45;
DFS[16'h0627] = 8'h86;
DFS[16'h0628] = 8'hC2;
DFS[16'h0629] = 8'h02;
DFS[16'h062A] = 8'hB0;
DFS[16'h062B] = 8'h26;
DFS[16'h062C] = 8'h00;
DFS[16'h062D] = 8'h42;
DFS[16'h062E] = 8'h55;
DFS[16'h062F] = 8'h49;
DFS[16'h0630] = 8'h4C;
DFS[16'h0631] = 8'h44;
DFS[16'h0632] = 8'h9F;
DFS[16'h0633] = 8'h47;
DFS[16'h0634] = 8'h01;
DFS[16'h0635] = 8'h43;
DFS[16'h0636] = 8'h41;
DFS[16'h0637] = 8'h52;
DFS[16'h0638] = 8'h44;
DFS[16'h0639] = 8'h93;
DFS[16'h063A] = 8'h37;
DFS[16'h063B] = 8'h00;
DFS[16'h063C] = 8'h44;
DFS[16'h063D] = 8'h55;
DFS[16'h063E] = 8'h4D;
DFS[16'h063F] = 8'h50;
DFS[16'h0640] = 8'h9E;
DFS[16'h0641] = 8'hCF;
DFS[16'h0642] = 8'h01;
DFS[16'h0643] = 8'h4C;
DFS[16'h0644] = 8'h49;
DFS[16'h0645] = 8'h53;
DFS[16'h0646] = 8'h54;
DFS[16'h0647] = 8'h9E;
DFS[16'h0648] = 8'h8D;
DFS[16'h0649] = 8'h01;
DFS[16'h064A] = 8'h54;
DFS[16'h064B] = 8'h59;
DFS[16'h064C] = 8'h50;
DFS[16'h064D] = 8'h45;
DFS[16'h064E] = 8'h9E;
DFS[16'h064F] = 8'h86;
DFS[16'h0650] = 8'h01;
DFS[16'h0651] = 8'h44;
DFS[16'h0652] = 8'h4D;
DFS[16'h0653] = 8'h4D;
DFS[16'h0654] = 8'h43;
DFS[16'h0655] = 8'h93;
DFS[16'h0656] = 8'h37;
DFS[16'h0657] = 8'h00;
DFS[16'h0658] = 8'h85;
DFS[16'h0659] = 8'hB6;
DFS[16'h065A] = 8'h00;
DFS[16'h065B] = 8'h44;
DFS[16'h065C] = 8'h46;
DFS[16'h065D] = 8'h53;
DFS[16'h065E] = 8'h99;
DFS[16'h065F] = 8'hC5;
DFS[16'h0660] = 8'h00;
DFS[16'h0661] = 8'h55;
DFS[16'h0662] = 8'h54;
DFS[16'h0663] = 8'h49;
DFS[16'h0664] = 8'h4C;
DFS[16'h0665] = 8'h53;
DFS[16'h0666] = 8'h99;
DFS[16'h0667] = 8'hED;
DFS[16'h0668] = 8'h00;
DFS[16'h0669] = 8'h99;
DFS[16'h066A] = 8'hF4;
DFS[16'h066B] = 8'h00;
DFS[16'h066C] = 8'h20;
DFS[16'h066D] = 8'hB8;
DFS[16'h066E] = 8'h86;
DFS[16'h066F] = 8'hA2;
DFS[16'h0670] = 8'hFD;
DFS[16'h0671] = 8'h8A;
DFS[16'h0672] = 8'hBA;
DFS[16'h0673] = 8'h86;
DFS[16'h0674] = 8'hB6;
DFS[16'h0675] = 8'hAA;
DFS[16'h0676] = 8'h98;
DFS[16'h0677] = 8'h48;
DFS[16'h0678] = 8'hE8;
DFS[16'h0679] = 8'hE8;
DFS[16'h067A] = 8'h68;
DFS[16'h067B] = 8'h48;
DFS[16'h067C] = 8'hA8;
DFS[16'h067D] = 8'h20;
DFS[16'h067E] = 8'hBF;
DFS[16'h067F] = 8'h86;
DFS[16'h0680] = 8'hE8;
DFS[16'h0681] = 8'hBD;
DFS[16'h0682] = 8'hB8;
DFS[16'h0683] = 8'h85;
DFS[16'h0684] = 8'h30;
DFS[16'h0685] = 8'h28;
DFS[16'h0686] = 8'hCA;
DFS[16'h0687] = 8'h88;
DFS[16'h0688] = 8'h86;
DFS[16'h0689] = 8'hB8;
DFS[16'h068A] = 8'hE8;
DFS[16'h068B] = 8'hC8;
DFS[16'h068C] = 8'hBD;
DFS[16'h068D] = 8'hB8;
DFS[16'h068E] = 8'h85;
DFS[16'h068F] = 8'h30;
DFS[16'h0690] = 8'h16;
DFS[16'h0691] = 8'h51;
DFS[16'h0692] = 8'hF2;
DFS[16'h0693] = 8'h29;
DFS[16'h0694] = 8'h5F;
DFS[16'h0695] = 8'hF0;
DFS[16'h0696] = 8'hF3;
DFS[16'h0697] = 8'hCA;
DFS[16'h0698] = 8'hE8;
DFS[16'h0699] = 8'hBD;
DFS[16'h069A] = 8'hB8;
DFS[16'h069B] = 8'h85;
DFS[16'h069C] = 8'h10;
DFS[16'h069D] = 8'hFA;
DFS[16'h069E] = 8'hB1;
DFS[16'h069F] = 8'hF2;
DFS[16'h06A0] = 8'hC9;
DFS[16'h06A1] = 8'h2E;
DFS[16'h06A2] = 8'hD0;
DFS[16'h06A3] = 8'hD4;
DFS[16'h06A4] = 8'hC8;
DFS[16'h06A5] = 8'hB0;
DFS[16'h06A6] = 8'h07;
DFS[16'h06A7] = 8'hB1;
DFS[16'h06A8] = 8'hF2;
DFS[16'h06A9] = 8'h20;
DFS[16'h06AA] = 8'hEE;
DFS[16'h06AB] = 8'h82;
DFS[16'h06AC] = 8'h90;
DFS[16'h06AD] = 8'hCA;
DFS[16'h06AE] = 8'h68;
DFS[16'h06AF] = 8'hBD;
DFS[16'h06B0] = 8'hB8;
DFS[16'h06B1] = 8'h85;
DFS[16'h06B2] = 8'h48;
DFS[16'h06B3] = 8'hBD;
DFS[16'h06B4] = 8'hB9;
DFS[16'h06B5] = 8'h85;
DFS[16'h06B6] = 8'h48;
DFS[16'h06B7] = 8'h60;
DFS[16'h06B8] = 8'h86;
DFS[16'h06B9] = 8'hF2;
DFS[16'h06BA] = 8'h84;
DFS[16'h06BB] = 8'hF3;
DFS[16'h06BC] = 8'hA0;
DFS[16'h06BD] = 8'h00;
DFS[16'h06BE] = 8'h60;
DFS[16'h06BF] = 8'h18;
DFS[16'h06C0] = 8'h4C;
DFS[16'h06C1] = 8'hC2;
DFS[16'h06C2] = 8'hFF;
DFS[16'h06C3] = 8'h20;
DFS[16'h06C4] = 8'h5E;
DFS[16'h06C5] = 8'h82;
DFS[16'h06C6] = 8'h20;
DFS[16'h06C7] = 8'h01;
DFS[16'h06C8] = 8'h9A;
DFS[16'h06C9] = 8'h20;
DFS[16'h06CA] = 8'h68;
DFS[16'h06CB] = 8'h82;
DFS[16'h06CC] = 8'hB9;
DFS[16'h06CD] = 8'h0F;
DFS[16'h06CE] = 8'h0E;
DFS[16'h06CF] = 8'h30;
DFS[16'h06D0] = 8'h12;
DFS[16'h06D1] = 8'h20;
DFS[16'h06D2] = 8'hC0;
DFS[16'h06D3] = 8'h81;
DFS[16'h06D4] = 8'h20;
DFS[16'h06D5] = 8'h65;
DFS[16'h06D6] = 8'h80;
DFS[16'h06D7] = 8'h20;
DFS[16'h06D8] = 8'h3A;
DFS[16'h06D9] = 8'h20;
DFS[16'h06DA] = 8'hEA;
DFS[16'h06DB] = 8'h20;
DFS[16'h06DC] = 8'h9E;
DFS[16'h06DD] = 8'h9C;
DFS[16'h06DE] = 8'hF0;
DFS[16'h06DF] = 8'h09;
DFS[16'h06E0] = 8'h20;
DFS[16'h06E1] = 8'h9A;
DFS[16'h06E2] = 8'h9F;
DFS[16'h06E3] = 8'h20;
DFS[16'h06E4] = 8'h9D;
DFS[16'h06E5] = 8'h82;
DFS[16'h06E6] = 8'hB0;
DFS[16'h06E7] = 8'hE4;
DFS[16'h06E8] = 8'h60;
DFS[16'h06E9] = 8'h20;
DFS[16'h06EA] = 8'hA1;
DFS[16'h06EB] = 8'h81;
DFS[16'h06EC] = 8'h20;
DFS[16'h06ED] = 8'hD1;
DFS[16'h06EE] = 8'h82;
DFS[16'h06EF] = 8'h20;
DFS[16'h06F0] = 8'hB4;
DFS[16'h06F1] = 8'h8A;
DFS[16'h06F2] = 8'hAC;
DFS[16'h06F3] = 8'hCE;
DFS[16'h06F4] = 8'h10;
DFS[16'h06F5] = 8'h20;
DFS[16'h06F6] = 8'h19;
DFS[16'h06F7] = 8'h82;
DFS[16'h06F8] = 8'h8C;
DFS[16'h06F9] = 8'hCE;
DFS[16'h06FA] = 8'h10;
DFS[16'h06FB] = 8'h4C;
DFS[16'h06FC] = 8'hE0;
DFS[16'h06FD] = 8'h86;
DFS[16'h06FE] = 8'h20;
DFS[16'h06FF] = 8'h62;
DFS[16'h0700] = 8'h82;
DFS[16'h0701] = 8'h20;
DFS[16'h0702] = 8'h01;
DFS[16'h0703] = 8'h9A;
DFS[16'h0704] = 8'h20;
DFS[16'h0705] = 8'h68;
DFS[16'h0706] = 8'h82;
DFS[16'h0707] = 8'h20;
DFS[16'h0708] = 8'hFC;
DFS[16'h0709] = 8'h82;
DFS[16'h070A] = 8'h20;
DFS[16'h070B] = 8'hD1;
DFS[16'h070C] = 8'h82;
DFS[16'h070D] = 8'h4C;
DFS[16'h070E] = 8'hB4;
DFS[16'h070F] = 8'h8A;
DFS[16'h0710] = 8'h20;
DFS[16'h0711] = 8'hBD;
DFS[16'h0712] = 8'h9B;
DFS[16'h0713] = 8'h20;
DFS[16'h0714] = 8'h5E;
DFS[16'h0715] = 8'h82;
DFS[16'h0716] = 8'h20;
DFS[16'h0717] = 8'h01;
DFS[16'h0718] = 8'h9A;
DFS[16'h0719] = 8'h20;
DFS[16'h071A] = 8'h68;
DFS[16'h071B] = 8'h82;
DFS[16'h071C] = 8'hB9;
DFS[16'h071D] = 8'h0F;
DFS[16'h071E] = 8'h0E;
DFS[16'h071F] = 8'h30;
DFS[16'h0720] = 8'h06;
DFS[16'h0721] = 8'h20;
DFS[16'h0722] = 8'hC0;
DFS[16'h0723] = 8'h81;
DFS[16'h0724] = 8'h20;
DFS[16'h0725] = 8'h9A;
DFS[16'h0726] = 8'h9F;
DFS[16'h0727] = 8'h20;
DFS[16'h0728] = 8'h9D;
DFS[16'h0729] = 8'h82;
DFS[16'h072A] = 8'hB0;
DFS[16'h072B] = 8'hF0;
DFS[16'h072C] = 8'h20;
DFS[16'h072D] = 8'h65;
DFS[16'h072E] = 8'h80;
DFS[16'h072F] = 8'h0D;
DFS[16'h0730] = 8'h44;
DFS[16'h0731] = 8'h65;
DFS[16'h0732] = 8'h6C;
DFS[16'h0733] = 8'h65;
DFS[16'h0734] = 8'h74;
DFS[16'h0735] = 8'h65;
DFS[16'h0736] = 8'h20;
DFS[16'h0737] = 8'h28;
DFS[16'h0738] = 8'h59;
DFS[16'h0739] = 8'h2F;
DFS[16'h073A] = 8'h4E;
DFS[16'h073B] = 8'h29;
DFS[16'h073C] = 8'h20;
DFS[16'h073D] = 8'h3F;
DFS[16'h073E] = 8'h20;
DFS[16'h073F] = 8'hEA;
DFS[16'h0740] = 8'h20;
DFS[16'h0741] = 8'h9E;
DFS[16'h0742] = 8'h9C;
DFS[16'h0743] = 8'hF0;
DFS[16'h0744] = 8'h03;
DFS[16'h0745] = 8'h4C;
DFS[16'h0746] = 8'h9A;
DFS[16'h0747] = 8'h9F;
DFS[16'h0748] = 8'h20;
DFS[16'h0749] = 8'hA1;
DFS[16'h074A] = 8'h81;
DFS[16'h074B] = 8'h20;
DFS[16'h074C] = 8'h96;
DFS[16'h074D] = 8'h82;
DFS[16'h074E] = 8'hB9;
DFS[16'h074F] = 8'h0F;
DFS[16'h0750] = 8'h0E;
DFS[16'h0751] = 8'h30;
DFS[16'h0752] = 8'h0C;
DFS[16'h0753] = 8'h20;
DFS[16'h0754] = 8'hD1;
DFS[16'h0755] = 8'h82;
DFS[16'h0756] = 8'hAC;
DFS[16'h0757] = 8'hCE;
DFS[16'h0758] = 8'h10;
DFS[16'h0759] = 8'h20;
DFS[16'h075A] = 8'h19;
DFS[16'h075B] = 8'h82;
DFS[16'h075C] = 8'h8C;
DFS[16'h075D] = 8'hCE;
DFS[16'h075E] = 8'h10;
DFS[16'h075F] = 8'h20;
DFS[16'h0760] = 8'h9D;
DFS[16'h0761] = 8'h82;
DFS[16'h0762] = 8'hB0;
DFS[16'h0763] = 8'hEA;
DFS[16'h0764] = 8'h20;
DFS[16'h0765] = 8'hB4;
DFS[16'h0766] = 8'h8A;
DFS[16'h0767] = 8'h20;
DFS[16'h0768] = 8'h65;
DFS[16'h0769] = 8'h80;
DFS[16'h076A] = 8'h0D;
DFS[16'h076B] = 8'h44;
DFS[16'h076C] = 8'h65;
DFS[16'h076D] = 8'h6C;
DFS[16'h076E] = 8'h65;
DFS[16'h076F] = 8'h74;
DFS[16'h0770] = 8'h65;
DFS[16'h0771] = 8'h64;
DFS[16'h0772] = 8'h0D;
DFS[16'h0773] = 8'hEA;
DFS[16'h0774] = 8'h60;
DFS[16'h0775] = 8'h20;
DFS[16'h0776] = 8'h01;
DFS[16'h0777] = 8'h9A;
DFS[16'h0778] = 8'h20;
DFS[16'h0779] = 8'h5D;
DFS[16'h077A] = 8'h83;
DFS[16'h077B] = 8'h8D;
DFS[16'h077C] = 8'hCB;
DFS[16'h077D] = 8'h10;
DFS[16'h077E] = 8'hEA;
DFS[16'h077F] = 8'hEA;
DFS[16'h0780] = 8'hEA;
DFS[16'h0781] = 8'h29;
DFS[16'h0782] = 8'h03;
DFS[16'h0783] = 8'h85;
DFS[16'h0784] = 8'hCF;
DFS[16'h0785] = 8'h60;
DFS[16'h0786] = 8'h20;
DFS[16'h0787] = 8'h61;
DFS[16'h0788] = 8'h89;
DFS[16'h0789] = 8'h20;
DFS[16'h078A] = 8'h6E;
DFS[16'h078B] = 8'h98;
DFS[16'h078C] = 8'h20;
DFS[16'h078D] = 8'h7E;
DFS[16'h078E] = 8'h83;
DFS[16'h078F] = 8'h4C;
DFS[16'h0790] = 8'hA5;
DFS[16'h0791] = 8'hAB;
DFS[16'h0792] = 8'hEA;
DFS[16'h0793] = 8'hEA;
DFS[16'h0794] = 8'h20;
DFS[16'h0795] = 8'h6E;
DFS[16'h0796] = 8'h82;
DFS[16'h0797] = 8'h20;
DFS[16'h0798] = 8'h6E;
DFS[16'h0799] = 8'h98;
DFS[16'h079A] = 8'h20;
DFS[16'h079B] = 8'h7E;
DFS[16'h079C] = 8'h83;
DFS[16'h079D] = 8'h84;
DFS[16'h079E] = 8'hBC;
DFS[16'h079F] = 8'hA2;
DFS[16'h07A0] = 8'h00;
DFS[16'h07A1] = 8'hA5;
DFS[16'h07A2] = 8'hC0;
DFS[16'h07A3] = 8'hD0;
DFS[16'h07A4] = 8'h06;
DFS[16'h07A5] = 8'hC8;
DFS[16'h07A6] = 8'hC8;
DFS[16'h07A7] = 8'hA2;
DFS[16'h07A8] = 8'h02;
DFS[16'h07A9] = 8'hD0;
DFS[16'h07AA] = 8'h08;
DFS[16'h07AB] = 8'hB9;
DFS[16'h07AC] = 8'h0E;
DFS[16'h07AD] = 8'h0F;
DFS[16'h07AE] = 8'h85;
DFS[16'h07AF] = 8'hC4;
DFS[16'h07B0] = 8'h20;
DFS[16'h07B1] = 8'h3F;
DFS[16'h07B2] = 8'h8A;
DFS[16'h07B3] = 8'hB9;
DFS[16'h07B4] = 8'h08;
DFS[16'h07B5] = 8'h0F;
DFS[16'h07B6] = 8'h95;
DFS[16'h07B7] = 8'hBE;
DFS[16'h07B8] = 8'hC8;
DFS[16'h07B9] = 8'hE8;
DFS[16'h07BA] = 8'hE0;
DFS[16'h07BB] = 8'h08;
DFS[16'h07BC] = 8'hD0;
DFS[16'h07BD] = 8'hF5;
DFS[16'h07BE] = 8'h20;
DFS[16'h07BF] = 8'h56;
DFS[16'h07C0] = 8'h8A;
DFS[16'h07C1] = 8'hA4;
DFS[16'h07C2] = 8'hBC;
DFS[16'h07C3] = 8'h20;
DFS[16'h07C4] = 8'hFC;
DFS[16'h07C5] = 8'h82;
DFS[16'h07C6] = 8'h4C;
DFS[16'h07C7] = 8'h96;
DFS[16'h07C8] = 8'hAB;
DFS[16'h07C9] = 8'h00;
DFS[16'h07CA] = 8'h00;
DFS[16'h07CB] = 8'h00;
DFS[16'h07CC] = 8'h00;
DFS[16'h07CD] = 8'h00;
DFS[16'h07CE] = 8'h00;
DFS[16'h07CF] = 8'h00;
DFS[16'h07D0] = 8'h00;
DFS[16'h07D1] = 8'h00;
DFS[16'h07D2] = 8'h00;
DFS[16'h07D3] = 8'h00;
DFS[16'h07D4] = 8'h20;
DFS[16'h07D5] = 8'hB8;
DFS[16'h07D6] = 8'h86;
DFS[16'h07D7] = 8'h20;
DFS[16'h07D8] = 8'h41;
DFS[16'h07D9] = 8'h88;
DFS[16'h07DA] = 8'h8C;
DFS[16'h07DB] = 8'hDB;
DFS[16'h07DC] = 8'h10;
DFS[16'h07DD] = 8'h20;
DFS[16'h07DE] = 8'h06;
DFS[16'h07DF] = 8'h81;
DFS[16'h07E0] = 8'h8C;
DFS[16'h07E1] = 8'hDA;
DFS[16'h07E2] = 8'h10;
DFS[16'h07E3] = 8'h20;
DFS[16'h07E4] = 8'h96;
DFS[16'h07E5] = 8'h82;
DFS[16'h07E6] = 8'hB0;
DFS[16'h07E7] = 8'h22;
DFS[16'h07E8] = 8'hAC;
DFS[16'h07E9] = 8'hDB;
DFS[16'h07EA] = 8'h10;
DFS[16'h07EB] = 8'hAD;
DFS[16'h07EC] = 8'hCC;
DFS[16'h07ED] = 8'h10;
DFS[16'h07EE] = 8'h85;
DFS[16'h07EF] = 8'hCE;
DFS[16'h07F0] = 8'hAD;
DFS[16'h07F1] = 8'hCD;
DFS[16'h07F2] = 8'h10;
DFS[16'h07F3] = 8'h20;
DFS[16'h07F4] = 8'h7E;
DFS[16'h07F5] = 8'h87;
DFS[16'h07F6] = 8'h20;
DFS[16'h07F7] = 8'h09;
DFS[16'h07F8] = 8'h81;
DFS[16'h07F9] = 8'h20;
DFS[16'h07FA] = 8'h96;
DFS[16'h07FB] = 8'h82;
DFS[16'h07FC] = 8'hB0;
DFS[16'h07FD] = 8'h0C;
DFS[16'h07FE] = 8'h20;
DFS[16'h07FF] = 8'h22;
DFS[16'h0800] = 8'h80;
DFS[16'h0801] = 8'hFE;
DFS[16'h0802] = 8'h63;
DFS[16'h0803] = 8'h6F;
DFS[16'h0804] = 8'h6D;
DFS[16'h0805] = 8'h6D;
DFS[16'h0806] = 8'h61;
DFS[16'h0807] = 8'h6E;
DFS[16'h0808] = 8'h64;
DFS[16'h0809] = 8'h00;
DFS[16'h080A] = 8'h20;
DFS[16'h080B] = 8'h9D;
DFS[16'h080C] = 8'h87;
DFS[16'h080D] = 8'h18;
DFS[16'h080E] = 8'hAD;
DFS[16'h080F] = 8'hDA;
DFS[16'h0810] = 8'h10;
DFS[16'h0811] = 8'hA8;
DFS[16'h0812] = 8'h65;
DFS[16'h0813] = 8'hF2;
DFS[16'h0814] = 8'h8D;
DFS[16'h0815] = 8'hDA;
DFS[16'h0816] = 8'h10;
DFS[16'h0817] = 8'hA5;
DFS[16'h0818] = 8'hF3;
DFS[16'h0819] = 8'h69;
DFS[16'h081A] = 8'h00;
DFS[16'h081B] = 8'h8D;
DFS[16'h081C] = 8'hDB;
DFS[16'h081D] = 8'h10;
DFS[16'h081E] = 8'hAD;
DFS[16'h081F] = 8'h76;
DFS[16'h0820] = 8'h10;
DFS[16'h0821] = 8'h2D;
DFS[16'h0822] = 8'h77;
DFS[16'h0823] = 8'h10;
DFS[16'h0824] = 8'h0D;
DFS[16'h0825] = 8'hD7;
DFS[16'h0826] = 8'h10;
DFS[16'h0827] = 8'hC9;
DFS[16'h0828] = 8'hFF;
DFS[16'h0829] = 8'hF0;
DFS[16'h082A] = 8'h13;
DFS[16'h082B] = 8'hA5;
DFS[16'h082C] = 8'hC0;
DFS[16'h082D] = 8'h8D;
DFS[16'h082E] = 8'h74;
DFS[16'h082F] = 8'h10;
DFS[16'h0830] = 8'hA5;
DFS[16'h0831] = 8'hC1;
DFS[16'h0832] = 8'h8D;
DFS[16'h0833] = 8'h75;
DFS[16'h0834] = 8'h10;
DFS[16'h0835] = 8'hA2;
DFS[16'h0836] = 8'h74;
DFS[16'h0837] = 8'hA0;
DFS[16'h0838] = 8'h10;
DFS[16'h0839] = 8'hA9;
DFS[16'h083A] = 8'h04;
DFS[16'h083B] = 8'h4C;
DFS[16'h083C] = 8'h06;
DFS[16'h083D] = 8'h04;
DFS[16'h083E] = 8'h6C;
DFS[16'h083F] = 8'hC0;
DFS[16'h0840] = 8'h00;
DFS[16'h0841] = 8'hA9;
DFS[16'h0842] = 8'hFF;
DFS[16'h0843] = 8'h85;
DFS[16'h0844] = 8'hC0;
DFS[16'h0845] = 8'hA5;
DFS[16'h0846] = 8'hF2;
DFS[16'h0847] = 8'h85;
DFS[16'h0848] = 8'hBC;
DFS[16'h0849] = 8'hA5;
DFS[16'h084A] = 8'hF3;
DFS[16'h084B] = 8'h85;
DFS[16'h084C] = 8'hBD;
DFS[16'h084D] = 8'h60;
DFS[16'h084E] = 8'hA2;
DFS[16'h084F] = 8'h00;
DFS[16'h0850] = 8'hF0;
DFS[16'h0851] = 8'h02;
DFS[16'h0852] = 8'hA2;
DFS[16'h0853] = 8'h02;
DFS[16'h0854] = 8'h20;
DFS[16'h0855] = 8'h60;
DFS[16'h0856] = 8'h88;
DFS[16'h0857] = 8'h9D;
DFS[16'h0858] = 8'hCB;
DFS[16'h0859] = 8'h10;
DFS[16'h085A] = 8'hA5;
DFS[16'h085B] = 8'hCE;
DFS[16'h085C] = 8'h9D;
DFS[16'h085D] = 8'hCA;
DFS[16'h085E] = 8'h10;
DFS[16'h085F] = 8'h60;
DFS[16'h0860] = 8'hA9;
DFS[16'h0861] = 8'h24;
DFS[16'h0862] = 8'h85;
DFS[16'h0863] = 8'hCE;
DFS[16'h0864] = 8'h20;
DFS[16'h0865] = 8'hBF;
DFS[16'h0866] = 8'h86;
DFS[16'h0867] = 8'hD0;
DFS[16'h0868] = 8'h07;
DFS[16'h0869] = 8'hA9;
DFS[16'h086A] = 8'h00;
DFS[16'h086B] = 8'h20;
DFS[16'h086C] = 8'h7E;
DFS[16'h086D] = 8'h87;
DFS[16'h086E] = 8'hF0;
DFS[16'h086F] = 8'h30;
DFS[16'h0870] = 8'hAD;
DFS[16'h0871] = 8'hCB;
DFS[16'h0872] = 8'h10;
DFS[16'h0873] = 8'h20;
DFS[16'h0874] = 8'h7E;
DFS[16'h0875] = 8'h87;
DFS[16'h0876] = 8'h20;
DFS[16'h0877] = 8'hC5;
DFS[16'h0878] = 8'hFF;
DFS[16'h0879] = 8'hB0;
DFS[16'h087A] = 8'h10;
DFS[16'h087B] = 8'hC9;
DFS[16'h087C] = 8'h3A;
DFS[16'h087D] = 8'hD0;
DFS[16'h087E] = 8'h1A;
DFS[16'h087F] = 8'h20;
DFS[16'h0880] = 8'h5D;
DFS[16'h0881] = 8'h83;
DFS[16'h0882] = 8'h20;
DFS[16'h0883] = 8'hC5;
DFS[16'h0884] = 8'hFF;
DFS[16'h0885] = 8'hB0;
DFS[16'h0886] = 8'h19;
DFS[16'h0887] = 8'hC9;
DFS[16'h0888] = 8'h2E;
DFS[16'h0889] = 8'hF0;
DFS[16'h088A] = 8'hEB;
DFS[16'h088B] = 8'h20;
DFS[16'h088C] = 8'h22;
DFS[16'h088D] = 8'h80;
DFS[16'h088E] = 8'hCE;
DFS[16'h088F] = 8'h64;
DFS[16'h0890] = 8'h69;
DFS[16'h0891] = 8'h72;
DFS[16'h0892] = 8'h65;
DFS[16'h0893] = 8'h63;
DFS[16'h0894] = 8'h74;
DFS[16'h0895] = 8'h6F;
DFS[16'h0896] = 8'h72;
DFS[16'h0897] = 8'h79;
DFS[16'h0898] = 8'h00;
DFS[16'h0899] = 8'h85;
DFS[16'h089A] = 8'hCE;
DFS[16'h089B] = 8'h20;
DFS[16'h089C] = 8'hC5;
DFS[16'h089D] = 8'hFF;
DFS[16'h089E] = 8'h90;
DFS[16'h089F] = 8'hEB;
DFS[16'h08A0] = 8'hA5;
DFS[16'h08A1] = 8'hCF;
DFS[16'h08A2] = 8'h60;
DFS[16'h08A3] = 8'h20;
DFS[16'h08A4] = 8'h01;
DFS[16'h08A5] = 8'h9A;
DFS[16'h08A6] = 8'h20;
DFS[16'h08A7] = 8'h4D;
DFS[16'h08A8] = 8'h83;
DFS[16'h08A9] = 8'h20;
DFS[16'h08AA] = 8'h47;
DFS[16'h08AB] = 8'h83;
DFS[16'h08AC] = 8'h4C;
DFS[16'h08AD] = 8'hA7;
DFS[16'h08AE] = 8'hAE;
DFS[16'h08AF] = 8'h00;
DFS[16'h08B0] = 8'h20;
DFS[16'h08B1] = 8'hC6;
DFS[16'h08B2] = 8'h88;
DFS[16'h08B3] = 8'hCA;
DFS[16'h08B4] = 8'h10;
DFS[16'h08B5] = 8'hFA;
DFS[16'h08B6] = 8'hE8;
DFS[16'h08B7] = 8'h20;
DFS[16'h08B8] = 8'hC5;
DFS[16'h08B9] = 8'hFF;
DFS[16'h08BA] = 8'hB0;
DFS[16'h08BB] = 8'h07;
DFS[16'h08BC] = 8'h20;
DFS[16'h08BD] = 8'hC6;
DFS[16'h08BE] = 8'h88;
DFS[16'h08BF] = 8'hE0;
DFS[16'h08C0] = 8'h0B;
DFS[16'h08C1] = 8'h90;
DFS[16'h08C2] = 8'hF3;
DFS[16'h08C3] = 8'h4C;
DFS[16'h08C4] = 8'hB4;
DFS[16'h08C5] = 8'h8A;
DFS[16'h08C6] = 8'hE0;
DFS[16'h08C7] = 8'h08;
DFS[16'h08C8] = 8'h90;
DFS[16'h08C9] = 8'h04;
DFS[16'h08CA] = 8'h9D;
DFS[16'h08CB] = 8'hF8;
DFS[16'h08CC] = 8'h0E;
DFS[16'h08CD] = 8'h60;
DFS[16'h08CE] = 8'h9D;
DFS[16'h08CF] = 8'h00;
DFS[16'h08D0] = 8'h0E;
DFS[16'h08D1] = 8'h60;
DFS[16'h08D2] = 8'h20;
DFS[16'h08D3] = 8'h5E;
DFS[16'h08D4] = 8'h82;
DFS[16'h08D5] = 8'h20;
DFS[16'h08D6] = 8'h01;
DFS[16'h08D7] = 8'h9A;
DFS[16'h08D8] = 8'h20;
DFS[16'h08D9] = 8'hFE;
DFS[16'h08DA] = 8'h80;
DFS[16'h08DB] = 8'hA2;
DFS[16'h08DC] = 8'h00;
DFS[16'h08DD] = 8'h20;
DFS[16'h08DE] = 8'hBF;
DFS[16'h08DF] = 8'h86;
DFS[16'h08E0] = 8'hD0;
DFS[16'h08E1] = 8'h23;
DFS[16'h08E2] = 8'h86;
DFS[16'h08E3] = 8'hAA;
DFS[16'h08E4] = 8'h20;
DFS[16'h08E5] = 8'h96;
DFS[16'h08E6] = 8'h82;
DFS[16'h08E7] = 8'hB0;
DFS[16'h08E8] = 8'h03;
DFS[16'h08E9] = 8'h4C;
DFS[16'h08EA] = 8'h76;
DFS[16'h08EB] = 8'h82;
DFS[16'h08EC] = 8'h20;
DFS[16'h08ED] = 8'h4F;
DFS[16'h08EE] = 8'h98;
DFS[16'h08EF] = 8'hB9;
DFS[16'h08F0] = 8'h0F;
DFS[16'h08F1] = 8'h0E;
DFS[16'h08F2] = 8'h29;
DFS[16'h08F3] = 8'h7F;
DFS[16'h08F4] = 8'h05;
DFS[16'h08F5] = 8'hAA;
DFS[16'h08F6] = 8'h99;
DFS[16'h08F7] = 8'h0F;
DFS[16'h08F8] = 8'h0E;
DFS[16'h08F9] = 8'h20;
DFS[16'h08FA] = 8'hFC;
DFS[16'h08FB] = 8'h82;
DFS[16'h08FC] = 8'h20;
DFS[16'h08FD] = 8'h9D;
DFS[16'h08FE] = 8'h82;
DFS[16'h08FF] = 8'hB0;
DFS[16'h0900] = 8'hEB;
DFS[16'h0901] = 8'h90;
DFS[16'h0902] = 8'hC0;
DFS[16'h0903] = 8'hA2;
DFS[16'h0904] = 8'h80;
DFS[16'h0905] = 8'h20;
DFS[16'h0906] = 8'hC5;
DFS[16'h0907] = 8'hFF;
DFS[16'h0908] = 8'hB0;
DFS[16'h0909] = 8'hD8;
DFS[16'h090A] = 8'hC9;
DFS[16'h090B] = 8'h4C;
DFS[16'h090C] = 8'hF0;
DFS[16'h090D] = 8'hF5;
DFS[16'h090E] = 8'h20;
DFS[16'h090F] = 8'h22;
DFS[16'h0910] = 8'h80;
DFS[16'h0911] = 8'hCF;
DFS[16'h0912] = 8'h61;
DFS[16'h0913] = 8'h74;
DFS[16'h0914] = 8'h74;
DFS[16'h0915] = 8'h72;
DFS[16'h0916] = 8'h69;
DFS[16'h0917] = 8'h62;
DFS[16'h0918] = 8'h75;
DFS[16'h0919] = 8'h74;
DFS[16'h091A] = 8'h65;
DFS[16'h091B] = 8'h00;
DFS[16'h091C] = 8'h20;
DFS[16'h091D] = 8'hE1;
DFS[16'h091E] = 8'h83;
DFS[16'h091F] = 8'h8A;
DFS[16'h0920] = 8'hC9;
DFS[16'h0921] = 8'h04;
DFS[16'h0922] = 8'hF0;
DFS[16'h0923] = 8'h1A;
DFS[16'h0924] = 8'hC9;
DFS[16'h0925] = 8'h02;
DFS[16'h0926] = 8'h90;
DFS[16'h0927] = 8'h0B;
DFS[16'h0928] = 8'h20;
DFS[16'h0929] = 8'h22;
DFS[16'h092A] = 8'h80;
DFS[16'h092B] = 8'hCB;
DFS[16'h092C] = 8'h6F;
DFS[16'h092D] = 8'h70;
DFS[16'h092E] = 8'h74;
DFS[16'h092F] = 8'h69;
DFS[16'h0930] = 8'h6F;
DFS[16'h0931] = 8'h6E;
DFS[16'h0932] = 8'h00;
DFS[16'h0933] = 8'hA2;
DFS[16'h0934] = 8'hFF;
DFS[16'h0935] = 8'h98;
DFS[16'h0936] = 8'hF0;
DFS[16'h0937] = 8'h02;
DFS[16'h0938] = 8'hA2;
DFS[16'h0939] = 8'h00;
DFS[16'h093A] = 8'h8E;
DFS[16'h093B] = 8'hC7;
DFS[16'h093C] = 8'h10;
DFS[16'h093D] = 8'h60;
DFS[16'h093E] = 8'h98;
DFS[16'h093F] = 8'h48;
DFS[16'h0940] = 8'h20;
DFS[16'h0941] = 8'h4D;
DFS[16'h0942] = 8'h83;
DFS[16'h0943] = 8'h20;
DFS[16'h0944] = 8'h4D;
DFS[16'h0945] = 8'hAB;
DFS[16'h0946] = 8'h68;
DFS[16'h0947] = 8'h20;
DFS[16'h0948] = 8'h0B;
DFS[16'h0949] = 8'h82;
DFS[16'h094A] = 8'h4D;
DFS[16'h094B] = 8'h06;
DFS[16'h094C] = 8'h0F;
DFS[16'h094D] = 8'h29;
DFS[16'h094E] = 8'h30;
DFS[16'h094F] = 8'h4D;
DFS[16'h0950] = 8'h06;
DFS[16'h0951] = 8'h0F;
DFS[16'h0952] = 8'h8D;
DFS[16'h0953] = 8'h06;
DFS[16'h0954] = 8'h0F;
DFS[16'h0955] = 8'h4C;
DFS[16'h0956] = 8'hB4;
DFS[16'h0957] = 8'h8A;
DFS[16'h0958] = 8'h20;
DFS[16'h0959] = 8'h18;
DFS[16'h095A] = 8'h80;
DFS[16'h095B] = 8'hC6;
DFS[16'h095C] = 8'h66;
DFS[16'h095D] = 8'h75;
DFS[16'h095E] = 8'h6C;
DFS[16'h095F] = 8'h6C;
DFS[16'h0960] = 8'h00;
DFS[16'h0961] = 8'h20;
DFS[16'h0962] = 8'h06;
DFS[16'h0963] = 8'h81;
DFS[16'h0964] = 8'h20;
DFS[16'h0965] = 8'h96;
DFS[16'h0966] = 8'h82;
DFS[16'h0967] = 8'h90;
DFS[16'h0968] = 8'h03;
DFS[16'h0969] = 8'h20;
DFS[16'h096A] = 8'hD1;
DFS[16'h096B] = 8'h82;
DFS[16'h096C] = 8'hA5;
DFS[16'h096D] = 8'hC2;
DFS[16'h096E] = 8'h48;
DFS[16'h096F] = 8'hA5;
DFS[16'h0970] = 8'hC3;
DFS[16'h0971] = 8'h48;
DFS[16'h0972] = 8'h38;
DFS[16'h0973] = 8'hA5;
DFS[16'h0974] = 8'hC4;
DFS[16'h0975] = 8'hE5;
DFS[16'h0976] = 8'hC2;
DFS[16'h0977] = 8'h85;
DFS[16'h0978] = 8'hC2;
DFS[16'h0979] = 8'hA5;
DFS[16'h097A] = 8'hC5;
DFS[16'h097B] = 8'hE5;
DFS[16'h097C] = 8'hC3;
DFS[16'h097D] = 8'h85;
DFS[16'h097E] = 8'hC3;
DFS[16'h097F] = 8'hAD;
DFS[16'h0980] = 8'h7A;
DFS[16'h0981] = 8'h10;
DFS[16'h0982] = 8'hED;
DFS[16'h0983] = 8'h78;
DFS[16'h0984] = 8'h10;
DFS[16'h0985] = 8'h85;
DFS[16'h0986] = 8'hC6;
DFS[16'h0987] = 8'h20;
DFS[16'h0988] = 8'h9D;
DFS[16'h0989] = 8'h89;
DFS[16'h098A] = 8'hAD;
DFS[16'h098B] = 8'h79;
DFS[16'h098C] = 8'h10;
DFS[16'h098D] = 8'h8D;
DFS[16'h098E] = 8'h75;
DFS[16'h098F] = 8'h10;
DFS[16'h0990] = 8'hAD;
DFS[16'h0991] = 8'h78;
DFS[16'h0992] = 8'h10;
DFS[16'h0993] = 8'h8D;
DFS[16'h0994] = 8'h74;
DFS[16'h0995] = 8'h10;
DFS[16'h0996] = 8'h68;
DFS[16'h0997] = 8'h85;
DFS[16'h0998] = 8'hBF;
DFS[16'h0999] = 8'h68;
DFS[16'h099A] = 8'h85;
DFS[16'h099B] = 8'hBE;
DFS[16'h099C] = 8'h60;
DFS[16'h099D] = 8'hA9;
DFS[16'h099E] = 8'h00;
DFS[16'h099F] = 8'h85;
DFS[16'h09A0] = 8'hC4;
DFS[16'h09A1] = 8'hA9;
DFS[16'h09A2] = 8'h02;
DFS[16'h09A3] = 8'h85;
DFS[16'h09A4] = 8'hC5;
DFS[16'h09A5] = 8'hAC;
DFS[16'h09A6] = 8'h05;
DFS[16'h09A7] = 8'h0F;
DFS[16'h09A8] = 8'hF0;
DFS[16'h09A9] = 8'h2D;
DFS[16'h09AA] = 8'hC0;
DFS[16'h09AB] = 8'hF8;
DFS[16'h09AC] = 8'hB0;
DFS[16'h09AD] = 8'h56;
DFS[16'h09AE] = 8'h20;
DFS[16'h09AF] = 8'h9E;
DFS[16'h09B0] = 8'h85;
DFS[16'h09B1] = 8'h4C;
DFS[16'h09B2] = 8'hBC;
DFS[16'h09B3] = 8'h89;
DFS[16'h09B4] = 8'hF0;
DFS[16'h09B5] = 8'hA2;
DFS[16'h09B6] = 8'h20;
DFS[16'h09B7] = 8'h19;
DFS[16'h09B8] = 8'h82;
DFS[16'h09B9] = 8'h20;
DFS[16'h09BA] = 8'h7F;
DFS[16'h09BB] = 8'h85;
DFS[16'h09BC] = 8'h98;
DFS[16'h09BD] = 8'h90;
DFS[16'h09BE] = 8'hF5;
DFS[16'h09BF] = 8'h84;
DFS[16'h09C0] = 8'hB0;
DFS[16'h09C1] = 8'hAC;
DFS[16'h09C2] = 8'h05;
DFS[16'h09C3] = 8'h0F;
DFS[16'h09C4] = 8'hC4;
DFS[16'h09C5] = 8'hB0;
DFS[16'h09C6] = 8'hF0;
DFS[16'h09C7] = 8'h0F;
DFS[16'h09C8] = 8'hB9;
DFS[16'h09C9] = 8'h07;
DFS[16'h09CA] = 8'h0E;
DFS[16'h09CB] = 8'h99;
DFS[16'h09CC] = 8'h0F;
DFS[16'h09CD] = 8'h0E;
DFS[16'h09CE] = 8'hB9;
DFS[16'h09CF] = 8'h07;
DFS[16'h09D0] = 8'h0F;
DFS[16'h09D1] = 8'h99;
DFS[16'h09D2] = 8'h0F;
DFS[16'h09D3] = 8'h0F;
DFS[16'h09D4] = 8'h88;
DFS[16'h09D5] = 8'hB0;
DFS[16'h09D6] = 8'hED;
DFS[16'h09D7] = 8'hA2;
DFS[16'h09D8] = 8'h00;
DFS[16'h09D9] = 8'h20;
DFS[16'h09DA] = 8'h17;
DFS[16'h09DB] = 8'h8A;
DFS[16'h09DC] = 8'hB5;
DFS[16'h09DD] = 8'hC7;
DFS[16'h09DE] = 8'h99;
DFS[16'h09DF] = 8'h08;
DFS[16'h09E0] = 8'h0E;
DFS[16'h09E1] = 8'hC8;
DFS[16'h09E2] = 8'hE8;
DFS[16'h09E3] = 8'hE0;
DFS[16'h09E4] = 8'h08;
DFS[16'h09E5] = 8'hD0;
DFS[16'h09E6] = 8'hF5;
DFS[16'h09E7] = 8'hB5;
DFS[16'h09E8] = 8'hBD;
DFS[16'h09E9] = 8'h88;
DFS[16'h09EA] = 8'h99;
DFS[16'h09EB] = 8'h08;
DFS[16'h09EC] = 8'h0F;
DFS[16'h09ED] = 8'hCA;
DFS[16'h09EE] = 8'hD0;
DFS[16'h09EF] = 8'hF7;
DFS[16'h09F0] = 8'h20;
DFS[16'h09F1] = 8'hFC;
DFS[16'h09F2] = 8'h82;
DFS[16'h09F3] = 8'h98;
DFS[16'h09F4] = 8'h48;
DFS[16'h09F5] = 8'hAC;
DFS[16'h09F6] = 8'h05;
DFS[16'h09F7] = 8'h0F;
DFS[16'h09F8] = 8'h20;
DFS[16'h09F9] = 8'h10;
DFS[16'h09FA] = 8'h82;
DFS[16'h09FB] = 8'h8C;
DFS[16'h09FC] = 8'h05;
DFS[16'h09FD] = 8'h0F;
DFS[16'h09FE] = 8'h20;
DFS[16'h09FF] = 8'hB4;
DFS[16'h0A00] = 8'h8A;
DFS[16'h0A01] = 8'h68;
DFS[16'h0A02] = 8'hA8;
DFS[16'h0A03] = 8'h60;
DFS[16'h0A04] = 8'h20;
DFS[16'h0A05] = 8'h33;
DFS[16'h0A06] = 8'h80;
DFS[16'h0A07] = 8'hBE;
DFS[16'h0A08] = 8'h43;
DFS[16'h0A09] = 8'h61;
DFS[16'h0A0A] = 8'h74;
DFS[16'h0A0B] = 8'h61;
DFS[16'h0A0C] = 8'h6C;
DFS[16'h0A0D] = 8'h6F;
DFS[16'h0A0E] = 8'h67;
DFS[16'h0A0F] = 8'h75;
DFS[16'h0A10] = 8'h65;
DFS[16'h0A11] = 8'h20;
DFS[16'h0A12] = 8'h66;
DFS[16'h0A13] = 8'h75;
DFS[16'h0A14] = 8'h6C;
DFS[16'h0A15] = 8'h6C;
DFS[16'h0A16] = 8'h00;
DFS[16'h0A17] = 8'hAD;
DFS[16'h0A18] = 8'h76;
DFS[16'h0A19] = 8'h10;
DFS[16'h0A1A] = 8'h29;
DFS[16'h0A1B] = 8'h03;
DFS[16'h0A1C] = 8'h0A;
DFS[16'h0A1D] = 8'h0A;
DFS[16'h0A1E] = 8'h45;
DFS[16'h0A1F] = 8'hC6;
DFS[16'h0A20] = 8'h29;
DFS[16'h0A21] = 8'hFC;
DFS[16'h0A22] = 8'h45;
DFS[16'h0A23] = 8'hC6;
DFS[16'h0A24] = 8'h0A;
DFS[16'h0A25] = 8'h0A;
DFS[16'h0A26] = 8'h4D;
DFS[16'h0A27] = 8'h74;
DFS[16'h0A28] = 8'h10;
DFS[16'h0A29] = 8'h29;
DFS[16'h0A2A] = 8'hFC;
DFS[16'h0A2B] = 8'h4D;
DFS[16'h0A2C] = 8'h74;
DFS[16'h0A2D] = 8'h10;
DFS[16'h0A2E] = 8'h0A;
DFS[16'h0A2F] = 8'h0A;
DFS[16'h0A30] = 8'h45;
DFS[16'h0A31] = 8'hC4;
DFS[16'h0A32] = 8'h29;
DFS[16'h0A33] = 8'hFC;
DFS[16'h0A34] = 8'h45;
DFS[16'h0A35] = 8'hC4;
DFS[16'h0A36] = 8'h85;
DFS[16'h0A37] = 8'hC4;
DFS[16'h0A38] = 8'h60;
DFS[16'h0A39] = 8'hA9;
DFS[16'h0A3A] = 8'h01;
DFS[16'h0A3B] = 8'h8D;
DFS[16'h0A3C] = 8'hC8;
DFS[16'h0A3D] = 8'h10;
DFS[16'h0A3E] = 8'h60;
DFS[16'h0A3F] = 8'hA9;
DFS[16'h0A40] = 8'h00;
DFS[16'h0A41] = 8'h8D;
DFS[16'h0A42] = 8'h75;
DFS[16'h0A43] = 8'h10;
DFS[16'h0A44] = 8'hA5;
DFS[16'h0A45] = 8'hC4;
DFS[16'h0A46] = 8'h20;
DFS[16'h0A47] = 8'hFF;
DFS[16'h0A48] = 8'h81;
DFS[16'h0A49] = 8'hC9;
DFS[16'h0A4A] = 8'h03;
DFS[16'h0A4B] = 8'hD0;
DFS[16'h0A4C] = 8'h05;
DFS[16'h0A4D] = 8'hA9;
DFS[16'h0A4E] = 8'hFF;
DFS[16'h0A4F] = 8'h8D;
DFS[16'h0A50] = 8'h75;
DFS[16'h0A51] = 8'h10;
DFS[16'h0A52] = 8'h8D;
DFS[16'h0A53] = 8'h74;
DFS[16'h0A54] = 8'h10;
DFS[16'h0A55] = 8'h60;
DFS[16'h0A56] = 8'hA9;
DFS[16'h0A57] = 8'h00;
DFS[16'h0A58] = 8'h8D;
DFS[16'h0A59] = 8'h77;
DFS[16'h0A5A] = 8'h10;
DFS[16'h0A5B] = 8'hA5;
DFS[16'h0A5C] = 8'hC4;
DFS[16'h0A5D] = 8'h20;
DFS[16'h0A5E] = 8'hFB;
DFS[16'h0A5F] = 8'h81;
DFS[16'h0A60] = 8'hC9;
DFS[16'h0A61] = 8'h03;
DFS[16'h0A62] = 8'hD0;
DFS[16'h0A63] = 8'h05;
DFS[16'h0A64] = 8'hA9;
DFS[16'h0A65] = 8'hFF;
DFS[16'h0A66] = 8'h8D;
DFS[16'h0A67] = 8'h77;
DFS[16'h0A68] = 8'h10;
DFS[16'h0A69] = 8'h8D;
DFS[16'h0A6A] = 8'h76;
DFS[16'h0A6B] = 8'h10;
DFS[16'h0A6C] = 8'h60;
DFS[16'h0A6D] = 8'h20;
DFS[16'h0A6E] = 8'h62;
DFS[16'h0A6F] = 8'h82;
DFS[16'h0A70] = 8'h20;
DFS[16'h0A71] = 8'hBF;
DFS[16'h0A72] = 8'h86;
DFS[16'h0A73] = 8'hD0;
DFS[16'h0A74] = 8'h03;
DFS[16'h0A75] = 8'h4C;
DFS[16'h0A76] = 8'h06;
DFS[16'h0A77] = 8'h9A;
DFS[16'h0A78] = 8'h20;
DFS[16'h0A79] = 8'hFE;
DFS[16'h0A7A] = 8'h80;
DFS[16'h0A7B] = 8'h98;
DFS[16'h0A7C] = 8'h48;
DFS[16'h0A7D] = 8'h20;
DFS[16'h0A7E] = 8'h96;
DFS[16'h0A7F] = 8'h82;
DFS[16'h0A80] = 8'hB0;
DFS[16'h0A81] = 8'h03;
DFS[16'h0A82] = 8'h4C;
DFS[16'h0A83] = 8'h76;
DFS[16'h0A84] = 8'h82;
DFS[16'h0A85] = 8'h20;
DFS[16'h0A86] = 8'h4C;
DFS[16'h0A87] = 8'h98;
DFS[16'h0A88] = 8'h84;
DFS[16'h0A89] = 8'hB3;
DFS[16'h0A8A] = 8'h68;
DFS[16'h0A8B] = 8'hA8;
DFS[16'h0A8C] = 8'h20;
DFS[16'h0A8D] = 8'hBF;
DFS[16'h0A8E] = 8'h86;
DFS[16'h0A8F] = 8'hF0;
DFS[16'h0A90] = 8'hE4;
DFS[16'h0A91] = 8'h20;
DFS[16'h0A92] = 8'hFE;
DFS[16'h0A93] = 8'h80;
DFS[16'h0A94] = 8'h20;
DFS[16'h0A95] = 8'h96;
DFS[16'h0A96] = 8'h82;
DFS[16'h0A97] = 8'h90;
DFS[16'h0A98] = 8'h0B;
DFS[16'h0A99] = 8'h20;
DFS[16'h0A9A] = 8'h2B;
DFS[16'h0A9B] = 8'h80;
DFS[16'h0A9C] = 8'hC4;
DFS[16'h0A9D] = 8'h65;
DFS[16'h0A9E] = 8'h78;
DFS[16'h0A9F] = 8'h69;
DFS[16'h0AA0] = 8'h73;
DFS[16'h0AA1] = 8'h74;
DFS[16'h0AA2] = 8'h73;
DFS[16'h0AA3] = 8'h00;
DFS[16'h0AA4] = 8'hA4;
DFS[16'h0AA5] = 8'hB3;
DFS[16'h0AA6] = 8'h20;
DFS[16'h0AA7] = 8'h10;
DFS[16'h0AA8] = 8'h82;
DFS[16'h0AA9] = 8'hA2;
DFS[16'h0AAA] = 8'h07;
DFS[16'h0AAB] = 8'hB5;
DFS[16'h0AAC] = 8'hC7;
DFS[16'h0AAD] = 8'h99;
DFS[16'h0AAE] = 8'h07;
DFS[16'h0AAF] = 8'h0E;
DFS[16'h0AB0] = 8'h88;
DFS[16'h0AB1] = 8'hCA;
DFS[16'h0AB2] = 8'h10;
DFS[16'h0AB3] = 8'hF7;
DFS[16'h0AB4] = 8'h18;
DFS[16'h0AB5] = 8'hF8;
DFS[16'h0AB6] = 8'hAD;
DFS[16'h0AB7] = 8'h04;
DFS[16'h0AB8] = 8'h0F;
DFS[16'h0AB9] = 8'h69;
DFS[16'h0ABA] = 8'h01;
DFS[16'h0ABB] = 8'hD8;
DFS[16'h0ABC] = 8'h8D;
DFS[16'h0ABD] = 8'h04;
DFS[16'h0ABE] = 8'h0F;
DFS[16'h0ABF] = 8'h4C;
DFS[16'h0AC0] = 8'h61;
DFS[16'h0AC1] = 8'hAB;
DFS[16'h0AC2] = 8'hA9;
DFS[16'h0AC3] = 8'hFF;
DFS[16'h0AC4] = 8'h20;
DFS[16'h0AC5] = 8'h9E;
DFS[16'h0AC6] = 8'h06;
DFS[16'h0AC7] = 8'hAD;
DFS[16'h0AC8] = 8'hE3;
DFS[16'h0AC9] = 8'hFE;
DFS[16'h0ACA] = 8'hA9;
DFS[16'h0ACB] = 8'h00;
DFS[16'h0ACC] = 8'h20;
DFS[16'h0ACD] = 8'h95;
DFS[16'h0ACE] = 8'h06;
DFS[16'h0ACF] = 8'hA8;
DFS[16'h0AD0] = 8'hB1;
DFS[16'h0AD1] = 8'hFD;
DFS[16'h0AD2] = 8'h20;
DFS[16'h0AD3] = 8'h95;
DFS[16'h0AD4] = 8'h06;
DFS[16'h0AD5] = 8'hC8;
DFS[16'h0AD6] = 8'hB1;
DFS[16'h0AD7] = 8'hFD;
DFS[16'h0AD8] = 8'h20;
DFS[16'h0AD9] = 8'h95;
DFS[16'h0ADA] = 8'h06;
DFS[16'h0ADB] = 8'hAA;
DFS[16'h0ADC] = 8'hD0;
DFS[16'h0ADD] = 8'hF7;
DFS[16'h0ADE] = 8'hA2;
DFS[16'h0ADF] = 8'hFF;
DFS[16'h0AE0] = 8'h9A;
DFS[16'h0AE1] = 8'h58;
DFS[16'h0AE2] = 8'h2C;
DFS[16'h0AE3] = 8'hE0;
DFS[16'h0AE4] = 8'hFE;
DFS[16'h0AE5] = 8'h10;
DFS[16'h0AE6] = 8'h06;
DFS[16'h0AE7] = 8'hAD;
DFS[16'h0AE8] = 8'hE1;
DFS[16'h0AE9] = 8'hFE;
DFS[16'h0AEA] = 8'h20;
DFS[16'h0AEB] = 8'hEE;
DFS[16'h0AEC] = 8'hFF;
DFS[16'h0AED] = 8'h2C;
DFS[16'h0AEE] = 8'hE2;
DFS[16'h0AEF] = 8'hFE;
DFS[16'h0AF0] = 8'h10;
DFS[16'h0AF1] = 8'hF0;
DFS[16'h0AF2] = 8'h2C;
DFS[16'h0AF3] = 8'hE0;
DFS[16'h0AF4] = 8'hFE;
DFS[16'h0AF5] = 8'h30;
DFS[16'h0AF6] = 8'hF0;
DFS[16'h0AF7] = 8'hAE;
DFS[16'h0AF8] = 8'hE3;
DFS[16'h0AF9] = 8'hFE;
DFS[16'h0AFA] = 8'h86;
DFS[16'h0AFB] = 8'h51;
DFS[16'h0AFC] = 8'h6C;
DFS[16'h0AFD] = 8'h00;
DFS[16'h0AFE] = 8'h05;
DFS[16'h0AFF] = 8'h00;
DFS[16'h0B00] = 8'h80;
DFS[16'h0B01] = 8'h00;
DFS[16'h0B02] = 8'h00;
DFS[16'h0B03] = 8'h4C;
DFS[16'h0B04] = 8'h84;
DFS[16'h0B05] = 8'h04;
DFS[16'h0B06] = 8'h4C;
DFS[16'h0B07] = 8'hA7;
DFS[16'h0B08] = 8'h06;
DFS[16'h0B09] = 8'hC9;
DFS[16'h0B0A] = 8'h80;
DFS[16'h0B0B] = 8'h90;
DFS[16'h0B0C] = 8'h2B;
DFS[16'h0B0D] = 8'hC9;
DFS[16'h0B0E] = 8'hC0;
DFS[16'h0B0F] = 8'hB0;
DFS[16'h0B10] = 8'h1A;
DFS[16'h0B11] = 8'h09;
DFS[16'h0B12] = 8'h40;
DFS[16'h0B13] = 8'hC5;
DFS[16'h0B14] = 8'h15;
DFS[16'h0B15] = 8'hD0;
DFS[16'h0B16] = 8'h20;
DFS[16'h0B17] = 8'h08;
DFS[16'h0B18] = 8'h78;
DFS[16'h0B19] = 8'hA9;
DFS[16'h0B1A] = 8'h05;
DFS[16'h0B1B] = 8'h20;
DFS[16'h0B1C] = 8'h9E;
DFS[16'h0B1D] = 8'h06;
DFS[16'h0B1E] = 8'hA5;
DFS[16'h0B1F] = 8'h15;
DFS[16'h0B20] = 8'h20;
DFS[16'h0B21] = 8'h9E;
DFS[16'h0B22] = 8'h06;
DFS[16'h0B23] = 8'h28;
DFS[16'h0B24] = 8'hA9;
DFS[16'h0B25] = 8'h80;
DFS[16'h0B26] = 8'h85;
DFS[16'h0B27] = 8'h15;
DFS[16'h0B28] = 8'h85;
DFS[16'h0B29] = 8'h14;
DFS[16'h0B2A] = 8'h60;
DFS[16'h0B2B] = 8'h06;
DFS[16'h0B2C] = 8'h14;
DFS[16'h0B2D] = 8'hB0;
DFS[16'h0B2E] = 8'h06;
DFS[16'h0B2F] = 8'hC5;
DFS[16'h0B30] = 8'h15;
DFS[16'h0B31] = 8'hF0;
DFS[16'h0B32] = 8'h04;
DFS[16'h0B33] = 8'h18;
DFS[16'h0B34] = 8'h60;
DFS[16'h0B35] = 8'h85;
DFS[16'h0B36] = 8'h15;
DFS[16'h0B37] = 8'h60;
DFS[16'h0B38] = 8'h08;
DFS[16'h0B39] = 8'h78;
DFS[16'h0B3A] = 8'h84;
DFS[16'h0B3B] = 8'h13;
DFS[16'h0B3C] = 8'h86;
DFS[16'h0B3D] = 8'h12;
DFS[16'h0B3E] = 8'h20;
DFS[16'h0B3F] = 8'h9E;
DFS[16'h0B40] = 8'h06;
DFS[16'h0B41] = 8'hAA;
DFS[16'h0B42] = 8'hA0;
DFS[16'h0B43] = 8'h03;
DFS[16'h0B44] = 8'hA5;
DFS[16'h0B45] = 8'h15;
DFS[16'h0B46] = 8'h20;
DFS[16'h0B47] = 8'h9E;
DFS[16'h0B48] = 8'h06;
DFS[16'h0B49] = 8'hB1;
DFS[16'h0B4A] = 8'h12;
DFS[16'h0B4B] = 8'h20;
DFS[16'h0B4C] = 8'h9E;
DFS[16'h0B4D] = 8'h06;
DFS[16'h0B4E] = 8'h88;
DFS[16'h0B4F] = 8'h10;
DFS[16'h0B50] = 8'hF8;
DFS[16'h0B51] = 8'hA0;
DFS[16'h0B52] = 8'h18;
DFS[16'h0B53] = 8'h8C;
DFS[16'h0B54] = 8'hE0;
DFS[16'h0B55] = 8'hFE;
DFS[16'h0B56] = 8'hBD;
DFS[16'h0B57] = 8'h18;
DFS[16'h0B58] = 8'h05;
DFS[16'h0B59] = 8'h8D;
DFS[16'h0B5A] = 8'hE0;
DFS[16'h0B5B] = 8'hFE;
DFS[16'h0B5C] = 8'h4A;
DFS[16'h0B5D] = 8'h4A;
DFS[16'h0B5E] = 8'h90;
DFS[16'h0B5F] = 8'h06;
DFS[16'h0B60] = 8'h2C;
DFS[16'h0B61] = 8'hE5;
DFS[16'h0B62] = 8'hFE;
DFS[16'h0B63] = 8'h2C;
DFS[16'h0B64] = 8'hE5;
DFS[16'h0B65] = 8'hFE;
DFS[16'h0B66] = 8'h20;
DFS[16'h0B67] = 8'h9E;
DFS[16'h0B68] = 8'h06;
DFS[16'h0B69] = 8'h2C;
DFS[16'h0B6A] = 8'hE6;
DFS[16'h0B6B] = 8'hFE;
DFS[16'h0B6C] = 8'h50;
DFS[16'h0B6D] = 8'hFB;
DFS[16'h0B6E] = 8'hB0;
DFS[16'h0B6F] = 8'h0D;
DFS[16'h0B70] = 8'hE0;
DFS[16'h0B71] = 8'h04;
DFS[16'h0B72] = 8'hD0;
DFS[16'h0B73] = 8'h11;
DFS[16'h0B74] = 8'h20;
DFS[16'h0B75] = 8'h14;
DFS[16'h0B76] = 8'h04;
DFS[16'h0B77] = 8'h20;
DFS[16'h0B78] = 8'h95;
DFS[16'h0B79] = 8'h06;
DFS[16'h0B7A] = 8'h4C;
DFS[16'h0B7B] = 8'h32;
DFS[16'h0B7C] = 8'h00;
DFS[16'h0B7D] = 8'h4A;
DFS[16'h0B7E] = 8'h90;
DFS[16'h0B7F] = 8'h05;
DFS[16'h0B80] = 8'hA0;
DFS[16'h0B81] = 8'h88;
DFS[16'h0B82] = 8'h8C;
DFS[16'h0B83] = 8'hE0;
DFS[16'h0B84] = 8'hFE;
DFS[16'h0B85] = 8'h28;
DFS[16'h0B86] = 8'h60;
DFS[16'h0B87] = 8'h58;
DFS[16'h0B88] = 8'hB0;
DFS[16'h0B89] = 8'h11;
DFS[16'h0B8A] = 8'hD0;
DFS[16'h0B8B] = 8'h03;
DFS[16'h0B8C] = 8'h4C;
DFS[16'h0B8D] = 8'h9C;
DFS[16'h0B8E] = 8'h05;
DFS[16'h0B8F] = 8'hA2;
DFS[16'h0B90] = 8'h00;
DFS[16'h0B91] = 8'hA0;
DFS[16'h0B92] = 8'hFF;
DFS[16'h0B93] = 8'hA9;
DFS[16'h0B94] = 8'hFD;
DFS[16'h0B95] = 8'h20;
DFS[16'h0B96] = 8'hF4;
DFS[16'h0B97] = 8'hFF;
DFS[16'h0B98] = 8'h8A;
DFS[16'h0B99] = 8'hF0;
DFS[16'h0B9A] = 8'hD9;
DFS[16'h0B9B] = 8'hA9;
DFS[16'h0B9C] = 8'hFF;
DFS[16'h0B9D] = 8'h20;
DFS[16'h0B9E] = 8'h06;
DFS[16'h0B9F] = 8'h04;
DFS[16'h0BA0] = 8'h90;
DFS[16'h0BA1] = 8'hF9;
DFS[16'h0BA2] = 8'h20;
DFS[16'h0BA3] = 8'hD2;
DFS[16'h0BA4] = 8'h04;
DFS[16'h0BA5] = 8'hA9;
DFS[16'h0BA6] = 8'h07;
DFS[16'h0BA7] = 8'h20;
DFS[16'h0BA8] = 8'hCB;
DFS[16'h0BA9] = 8'h04;
DFS[16'h0BAA] = 8'hA0;
DFS[16'h0BAB] = 8'h00;
DFS[16'h0BAC] = 8'h84;
DFS[16'h0BAD] = 8'h00;
DFS[16'h0BAE] = 8'hB1;
DFS[16'h0BAF] = 8'h00;
DFS[16'h0BB0] = 8'h8D;
DFS[16'h0BB1] = 8'hE5;
DFS[16'h0BB2] = 8'hFE;
DFS[16'h0BB3] = 8'hEA;
DFS[16'h0BB4] = 8'hEA;
DFS[16'h0BB5] = 8'hEA;
DFS[16'h0BB6] = 8'hC8;
DFS[16'h0BB7] = 8'hD0;
DFS[16'h0BB8] = 8'hF5;
DFS[16'h0BB9] = 8'hE6;
DFS[16'h0BBA] = 8'h54;
DFS[16'h0BBB] = 8'hD0;
DFS[16'h0BBC] = 8'h06;
DFS[16'h0BBD] = 8'hE6;
DFS[16'h0BBE] = 8'h55;
DFS[16'h0BBF] = 8'hD0;
DFS[16'h0BC0] = 8'h02;
DFS[16'h0BC1] = 8'hE6;
DFS[16'h0BC2] = 8'h56;
DFS[16'h0BC3] = 8'hE6;
DFS[16'h0BC4] = 8'h01;
DFS[16'h0BC5] = 8'h24;
DFS[16'h0BC6] = 8'h01;
DFS[16'h0BC7] = 8'h50;
DFS[16'h0BC8] = 8'hDC;
DFS[16'h0BC9] = 8'h20;
DFS[16'h0BCA] = 8'hD2;
DFS[16'h0BCB] = 8'h04;
DFS[16'h0BCC] = 8'hA9;
DFS[16'h0BCD] = 8'h04;
DFS[16'h0BCE] = 8'hA0;
DFS[16'h0BCF] = 8'h00;
DFS[16'h0BD0] = 8'hA2;
DFS[16'h0BD1] = 8'h53;
DFS[16'h0BD2] = 8'h4C;
DFS[16'h0BD3] = 8'h06;
DFS[16'h0BD4] = 8'h04;
DFS[16'h0BD5] = 8'hA9;
DFS[16'h0BD6] = 8'h80;
DFS[16'h0BD7] = 8'h85;
DFS[16'h0BD8] = 8'h54;
DFS[16'h0BD9] = 8'h85;
DFS[16'h0BDA] = 8'h01;
DFS[16'h0BDB] = 8'hA9;
DFS[16'h0BDC] = 8'h20;
DFS[16'h0BDD] = 8'h2D;
DFS[16'h0BDE] = 8'h06;
DFS[16'h0BDF] = 8'h80;
DFS[16'h0BE0] = 8'hA8;
DFS[16'h0BE1] = 8'h84;
DFS[16'h0BE2] = 8'h53;
DFS[16'h0BE3] = 8'hF0;
DFS[16'h0BE4] = 8'h19;
DFS[16'h0BE5] = 8'hAE;
DFS[16'h0BE6] = 8'h07;
DFS[16'h0BE7] = 8'h80;
DFS[16'h0BE8] = 8'hE8;
DFS[16'h0BE9] = 8'hBD;
DFS[16'h0BEA] = 8'h00;
DFS[16'h0BEB] = 8'h80;
DFS[16'h0BEC] = 8'hD0;
DFS[16'h0BED] = 8'hFA;
DFS[16'h0BEE] = 8'hBD;
DFS[16'h0BEF] = 8'h01;
DFS[16'h0BF0] = 8'h80;
DFS[16'h0BF1] = 8'h85;
DFS[16'h0BF2] = 8'h53;
DFS[16'h0BF3] = 8'hBD;
DFS[16'h0BF4] = 8'h02;
DFS[16'h0BF5] = 8'h80;
DFS[16'h0BF6] = 8'h85;
DFS[16'h0BF7] = 8'h54;
DFS[16'h0BF8] = 8'hBC;
DFS[16'h0BF9] = 8'h03;
DFS[16'h0BFA] = 8'h80;
DFS[16'h0BFB] = 8'hBD;
DFS[16'h0BFC] = 8'h04;
DFS[16'h0BFD] = 8'h80;
DFS[16'h0BFE] = 8'h85;
DFS[16'h0BFF] = 8'h56;
DFS[16'h0C00] = 8'h84;
DFS[16'h0C01] = 8'h55;
DFS[16'h0C02] = 8'h60;
DFS[16'h0C03] = 8'h37;
DFS[16'h0C04] = 8'h05;
DFS[16'h0C05] = 8'h96;
DFS[16'h0C06] = 8'h05;
DFS[16'h0C07] = 8'hF2;
DFS[16'h0C08] = 8'h05;
DFS[16'h0C09] = 8'h07;
DFS[16'h0C0A] = 8'h06;
DFS[16'h0C0B] = 8'h27;
DFS[16'h0C0C] = 8'h06;
DFS[16'h0C0D] = 8'h68;
DFS[16'h0C0E] = 8'h06;
DFS[16'h0C0F] = 8'h5E;
DFS[16'h0C10] = 8'h05;
DFS[16'h0C11] = 8'h2D;
DFS[16'h0C12] = 8'h05;
DFS[16'h0C13] = 8'h20;
DFS[16'h0C14] = 8'h05;
DFS[16'h0C15] = 8'h42;
DFS[16'h0C16] = 8'h05;
DFS[16'h0C17] = 8'hA9;
DFS[16'h0C18] = 8'h05;
DFS[16'h0C19] = 8'hD1;
DFS[16'h0C1A] = 8'h05;
DFS[16'h0C1B] = 8'h86;
DFS[16'h0C1C] = 8'h88;
DFS[16'h0C1D] = 8'h96;
DFS[16'h0C1E] = 8'h98;
DFS[16'h0C1F] = 8'h18;
DFS[16'h0C20] = 8'h18;
DFS[16'h0C21] = 8'h82;
DFS[16'h0C22] = 8'h18;
DFS[16'h0C23] = 8'h20;
DFS[16'h0C24] = 8'hC5;
DFS[16'h0C25] = 8'h06;
DFS[16'h0C26] = 8'hA8;
DFS[16'h0C27] = 8'h20;
DFS[16'h0C28] = 8'hC5;
DFS[16'h0C29] = 8'h06;
DFS[16'h0C2A] = 8'h20;
DFS[16'h0C2B] = 8'hD4;
DFS[16'h0C2C] = 8'hFF;
DFS[16'h0C2D] = 8'h4C;
DFS[16'h0C2E] = 8'h9C;
DFS[16'h0C2F] = 8'h05;
DFS[16'h0C30] = 8'h20;
DFS[16'h0C31] = 8'hC5;
DFS[16'h0C32] = 8'h06;
DFS[16'h0C33] = 8'hA8;
DFS[16'h0C34] = 8'h20;
DFS[16'h0C35] = 8'hD7;
DFS[16'h0C36] = 8'hFF;
DFS[16'h0C37] = 8'h4C;
DFS[16'h0C38] = 8'h3A;
DFS[16'h0C39] = 8'h05;
DFS[16'h0C3A] = 8'h20;
DFS[16'h0C3B] = 8'hE0;
DFS[16'h0C3C] = 8'hFF;
DFS[16'h0C3D] = 8'h6A;
DFS[16'h0C3E] = 8'h20;
DFS[16'h0C3F] = 8'h95;
DFS[16'h0C40] = 8'h06;
DFS[16'h0C41] = 8'h2A;
DFS[16'h0C42] = 8'h4C;
DFS[16'h0C43] = 8'h9E;
DFS[16'h0C44] = 8'h05;
DFS[16'h0C45] = 8'h20;
DFS[16'h0C46] = 8'hC5;
DFS[16'h0C47] = 8'h06;
DFS[16'h0C48] = 8'hF0;
DFS[16'h0C49] = 8'h0B;
DFS[16'h0C4A] = 8'h48;
DFS[16'h0C4B] = 8'h20;
DFS[16'h0C4C] = 8'h82;
DFS[16'h0C4D] = 8'h05;
DFS[16'h0C4E] = 8'h68;
DFS[16'h0C4F] = 8'h20;
DFS[16'h0C50] = 8'hCE;
DFS[16'h0C51] = 8'hFF;
DFS[16'h0C52] = 8'h4C;
DFS[16'h0C53] = 8'h9E;
DFS[16'h0C54] = 8'h05;
DFS[16'h0C55] = 8'h20;
DFS[16'h0C56] = 8'hC5;
DFS[16'h0C57] = 8'h06;
DFS[16'h0C58] = 8'hA8;
DFS[16'h0C59] = 8'hA9;
DFS[16'h0C5A] = 8'h00;
DFS[16'h0C5B] = 8'h20;
DFS[16'h0C5C] = 8'hCE;
DFS[16'h0C5D] = 8'hFF;
DFS[16'h0C5E] = 8'h4C;
DFS[16'h0C5F] = 8'h9C;
DFS[16'h0C60] = 8'h05;
DFS[16'h0C61] = 8'h20;
DFS[16'h0C62] = 8'hC5;
DFS[16'h0C63] = 8'h06;
DFS[16'h0C64] = 8'hA8;
DFS[16'h0C65] = 8'hA2;
DFS[16'h0C66] = 8'h04;
DFS[16'h0C67] = 8'h20;
DFS[16'h0C68] = 8'hC5;
DFS[16'h0C69] = 8'h06;
DFS[16'h0C6A] = 8'h95;
DFS[16'h0C6B] = 8'hFF;
DFS[16'h0C6C] = 8'hCA;
DFS[16'h0C6D] = 8'hD0;
DFS[16'h0C6E] = 8'hF8;
DFS[16'h0C6F] = 8'h20;
DFS[16'h0C70] = 8'hC5;
DFS[16'h0C71] = 8'h06;
DFS[16'h0C72] = 8'h20;
DFS[16'h0C73] = 8'hDA;
DFS[16'h0C74] = 8'hFF;
DFS[16'h0C75] = 8'h20;
DFS[16'h0C76] = 8'h95;
DFS[16'h0C77] = 8'h06;
DFS[16'h0C78] = 8'hA2;
DFS[16'h0C79] = 8'h03;
DFS[16'h0C7A] = 8'hB5;
DFS[16'h0C7B] = 8'h00;
DFS[16'h0C7C] = 8'h20;
DFS[16'h0C7D] = 8'h95;
DFS[16'h0C7E] = 8'h06;
DFS[16'h0C7F] = 8'hCA;
DFS[16'h0C80] = 8'h10;
DFS[16'h0C81] = 8'hF8;
DFS[16'h0C82] = 8'h4C;
DFS[16'h0C83] = 8'h36;
DFS[16'h0C84] = 8'h00;
DFS[16'h0C85] = 8'hA2;
DFS[16'h0C86] = 8'h00;
DFS[16'h0C87] = 8'hA0;
DFS[16'h0C88] = 8'h00;
DFS[16'h0C89] = 8'h20;
DFS[16'h0C8A] = 8'hC5;
DFS[16'h0C8B] = 8'h06;
DFS[16'h0C8C] = 8'h99;
DFS[16'h0C8D] = 8'h00;
DFS[16'h0C8E] = 8'h07;
DFS[16'h0C8F] = 8'hC8;
DFS[16'h0C90] = 8'hF0;
DFS[16'h0C91] = 8'h04;
DFS[16'h0C92] = 8'hC9;
DFS[16'h0C93] = 8'h0D;
DFS[16'h0C94] = 8'hD0;
DFS[16'h0C95] = 8'hF3;
DFS[16'h0C96] = 8'hA0;
DFS[16'h0C97] = 8'h07;
DFS[16'h0C98] = 8'h60;
DFS[16'h0C99] = 8'h20;
DFS[16'h0C9A] = 8'h82;
DFS[16'h0C9B] = 8'h05;
DFS[16'h0C9C] = 8'h20;
DFS[16'h0C9D] = 8'hF7;
DFS[16'h0C9E] = 8'hFF;
DFS[16'h0C9F] = 8'hA9;
DFS[16'h0CA0] = 8'h7F;
DFS[16'h0CA1] = 8'h2C;
DFS[16'h0CA2] = 8'hE2;
DFS[16'h0CA3] = 8'hFE;
DFS[16'h0CA4] = 8'h50;
DFS[16'h0CA5] = 8'hFB;
DFS[16'h0CA6] = 8'h8D;
DFS[16'h0CA7] = 8'hE3;
DFS[16'h0CA8] = 8'hFE;
DFS[16'h0CA9] = 8'h4C;
DFS[16'h0CAA] = 8'h36;
DFS[16'h0CAB] = 8'h00;
DFS[16'h0CAC] = 8'hA2;
DFS[16'h0CAD] = 8'h10;
DFS[16'h0CAE] = 8'h20;
DFS[16'h0CAF] = 8'hC5;
DFS[16'h0CB0] = 8'h06;
DFS[16'h0CB1] = 8'h95;
DFS[16'h0CB2] = 8'h01;
DFS[16'h0CB3] = 8'hCA;
DFS[16'h0CB4] = 8'hD0;
DFS[16'h0CB5] = 8'hF8;
DFS[16'h0CB6] = 8'h20;
DFS[16'h0CB7] = 8'h82;
DFS[16'h0CB8] = 8'h05;
DFS[16'h0CB9] = 8'h86;
DFS[16'h0CBA] = 8'h00;
DFS[16'h0CBB] = 8'h84;
DFS[16'h0CBC] = 8'h01;
DFS[16'h0CBD] = 8'hA0;
DFS[16'h0CBE] = 8'h00;
DFS[16'h0CBF] = 8'h20;
DFS[16'h0CC0] = 8'hC5;
DFS[16'h0CC1] = 8'h06;
DFS[16'h0CC2] = 8'h20;
DFS[16'h0CC3] = 8'hDD;
DFS[16'h0CC4] = 8'hFF;
DFS[16'h0CC5] = 8'h20;
DFS[16'h0CC6] = 8'h95;
DFS[16'h0CC7] = 8'h06;
DFS[16'h0CC8] = 8'hA2;
DFS[16'h0CC9] = 8'h10;
DFS[16'h0CCA] = 8'hB5;
DFS[16'h0CCB] = 8'h01;
DFS[16'h0CCC] = 8'h20;
DFS[16'h0CCD] = 8'h95;
DFS[16'h0CCE] = 8'h06;
DFS[16'h0CCF] = 8'hCA;
DFS[16'h0CD0] = 8'hD0;
DFS[16'h0CD1] = 8'hF8;
DFS[16'h0CD2] = 8'hF0;
DFS[16'h0CD3] = 8'hD5;
DFS[16'h0CD4] = 8'hA2;
DFS[16'h0CD5] = 8'h0D;
DFS[16'h0CD6] = 8'h20;
DFS[16'h0CD7] = 8'hC5;
DFS[16'h0CD8] = 8'h06;
DFS[16'h0CD9] = 8'h95;
DFS[16'h0CDA] = 8'hFF;
DFS[16'h0CDB] = 8'hCA;
DFS[16'h0CDC] = 8'hD0;
DFS[16'h0CDD] = 8'hF8;
DFS[16'h0CDE] = 8'h20;
DFS[16'h0CDF] = 8'hC5;
DFS[16'h0CE0] = 8'h06;
DFS[16'h0CE1] = 8'hA0;
DFS[16'h0CE2] = 8'h00;
DFS[16'h0CE3] = 8'h20;
DFS[16'h0CE4] = 8'hD1;
DFS[16'h0CE5] = 8'hFF;
DFS[16'h0CE6] = 8'h48;
DFS[16'h0CE7] = 8'hA2;
DFS[16'h0CE8] = 8'h0C;
DFS[16'h0CE9] = 8'hB5;
DFS[16'h0CEA] = 8'h00;
DFS[16'h0CEB] = 8'h20;
DFS[16'h0CEC] = 8'h95;
DFS[16'h0CED] = 8'h06;
DFS[16'h0CEE] = 8'hCA;
DFS[16'h0CEF] = 8'h10;
DFS[16'h0CF0] = 8'hF8;
DFS[16'h0CF1] = 8'h68;
DFS[16'h0CF2] = 8'h4C;
DFS[16'h0CF3] = 8'h3A;
DFS[16'h0CF4] = 8'h05;
DFS[16'h0CF5] = 8'h20;
DFS[16'h0CF6] = 8'hC5;
DFS[16'h0CF7] = 8'h06;
DFS[16'h0CF8] = 8'hAA;
DFS[16'h0CF9] = 8'h20;
DFS[16'h0CFA] = 8'hC5;
DFS[16'h0CFB] = 8'h06;
DFS[16'h0CFC] = 8'h20;
DFS[16'h0CFD] = 8'hF4;
DFS[16'h0CFE] = 8'hFF;
DFS[16'h0CFF] = 8'h2C;
DFS[16'h0D00] = 8'hE2;
DFS[16'h0D01] = 8'hFE;
DFS[16'h0D02] = 8'h50;
DFS[16'h0D03] = 8'hFB;
DFS[16'h0D04] = 8'h8E;
DFS[16'h0D05] = 8'hE3;
DFS[16'h0D06] = 8'hFE;
DFS[16'h0D07] = 8'h4C;
DFS[16'h0D08] = 8'h36;
DFS[16'h0D09] = 8'h00;
DFS[16'h0D0A] = 8'h20;
DFS[16'h0D0B] = 8'hC5;
DFS[16'h0D0C] = 8'h06;
DFS[16'h0D0D] = 8'hAA;
DFS[16'h0D0E] = 8'h20;
DFS[16'h0D0F] = 8'hC5;
DFS[16'h0D10] = 8'h06;
DFS[16'h0D11] = 8'hA8;
DFS[16'h0D12] = 8'h20;
DFS[16'h0D13] = 8'hC5;
DFS[16'h0D14] = 8'h06;
DFS[16'h0D15] = 8'h20;
DFS[16'h0D16] = 8'hF4;
DFS[16'h0D17] = 8'hFF;
DFS[16'h0D18] = 8'h49;
DFS[16'h0D19] = 8'h9D;
DFS[16'h0D1A] = 8'hF0;
DFS[16'h0D1B] = 8'hEB;
DFS[16'h0D1C] = 8'h6A;
DFS[16'h0D1D] = 8'h20;
DFS[16'h0D1E] = 8'h95;
DFS[16'h0D1F] = 8'h06;
DFS[16'h0D20] = 8'h2C;
DFS[16'h0D21] = 8'hE2;
DFS[16'h0D22] = 8'hFE;
DFS[16'h0D23] = 8'h50;
DFS[16'h0D24] = 8'hFB;
DFS[16'h0D25] = 8'h8C;
DFS[16'h0D26] = 8'hE3;
DFS[16'h0D27] = 8'hFE;
DFS[16'h0D28] = 8'h70;
DFS[16'h0D29] = 8'hD5;
DFS[16'h0D2A] = 8'h20;
DFS[16'h0D2B] = 8'hC5;
DFS[16'h0D2C] = 8'h06;
DFS[16'h0D2D] = 8'hA8;
DFS[16'h0D2E] = 8'h2C;
DFS[16'h0D2F] = 8'hE2;
DFS[16'h0D30] = 8'hFE;
DFS[16'h0D31] = 8'h10;
DFS[16'h0D32] = 8'hFB;
DFS[16'h0D33] = 8'hAE;
DFS[16'h0D34] = 8'hE3;
DFS[16'h0D35] = 8'hFE;
DFS[16'h0D36] = 8'hCA;
DFS[16'h0D37] = 8'h30;
DFS[16'h0D38] = 8'h0F;
DFS[16'h0D39] = 8'h2C;
DFS[16'h0D3A] = 8'hE2;
DFS[16'h0D3B] = 8'hFE;
DFS[16'h0D3C] = 8'h10;
DFS[16'h0D3D] = 8'hFB;
DFS[16'h0D3E] = 8'hAD;
DFS[16'h0D3F] = 8'hE3;
DFS[16'h0D40] = 8'hFE;
DFS[16'h0D41] = 8'h9D;
DFS[16'h0D42] = 8'h28;
DFS[16'h0D43] = 8'h01;
DFS[16'h0D44] = 8'hCA;
DFS[16'h0D45] = 8'h10;
DFS[16'h0D46] = 8'hF2;
DFS[16'h0D47] = 8'h98;
DFS[16'h0D48] = 8'hA2;
DFS[16'h0D49] = 8'h28;
DFS[16'h0D4A] = 8'hA0;
DFS[16'h0D4B] = 8'h01;
DFS[16'h0D4C] = 8'h20;
DFS[16'h0D4D] = 8'hF1;
DFS[16'h0D4E] = 8'hFF;
DFS[16'h0D4F] = 8'h2C;
DFS[16'h0D50] = 8'hE2;
DFS[16'h0D51] = 8'hFE;
DFS[16'h0D52] = 8'h10;
DFS[16'h0D53] = 8'hFB;
DFS[16'h0D54] = 8'hAE;
DFS[16'h0D55] = 8'hE3;
DFS[16'h0D56] = 8'hFE;
DFS[16'h0D57] = 8'hCA;
DFS[16'h0D58] = 8'h30;
DFS[16'h0D59] = 8'h0E;
DFS[16'h0D5A] = 8'hBC;
DFS[16'h0D5B] = 8'h28;
DFS[16'h0D5C] = 8'h01;
DFS[16'h0D5D] = 8'h2C;
DFS[16'h0D5E] = 8'hE2;
DFS[16'h0D5F] = 8'hFE;
DFS[16'h0D60] = 8'h50;
DFS[16'h0D61] = 8'hFB;
DFS[16'h0D62] = 8'h8C;
DFS[16'h0D63] = 8'hE3;
DFS[16'h0D64] = 8'hFE;
DFS[16'h0D65] = 8'hCA;
DFS[16'h0D66] = 8'h10;
DFS[16'h0D67] = 8'hF2;
DFS[16'h0D68] = 8'h4C;
DFS[16'h0D69] = 8'h36;
DFS[16'h0D6A] = 8'h00;
DFS[16'h0D6B] = 8'hA2;
DFS[16'h0D6C] = 8'h04;
DFS[16'h0D6D] = 8'h20;
DFS[16'h0D6E] = 8'hC5;
DFS[16'h0D6F] = 8'h06;
DFS[16'h0D70] = 8'h95;
DFS[16'h0D71] = 8'h00;
DFS[16'h0D72] = 8'hCA;
DFS[16'h0D73] = 8'h10;
DFS[16'h0D74] = 8'hF8;
DFS[16'h0D75] = 8'hE8;
DFS[16'h0D76] = 8'hA0;
DFS[16'h0D77] = 8'h00;
DFS[16'h0D78] = 8'h8A;
DFS[16'h0D79] = 8'h20;
DFS[16'h0D7A] = 8'hF1;
DFS[16'h0D7B] = 8'hFF;
DFS[16'h0D7C] = 8'h90;
DFS[16'h0D7D] = 8'h05;
DFS[16'h0D7E] = 8'hA9;
DFS[16'h0D7F] = 8'hFF;
DFS[16'h0D80] = 8'h4C;
DFS[16'h0D81] = 8'h9E;
DFS[16'h0D82] = 8'h05;
DFS[16'h0D83] = 8'hA2;
DFS[16'h0D84] = 8'h00;
DFS[16'h0D85] = 8'hA9;
DFS[16'h0D86] = 8'h7F;
DFS[16'h0D87] = 8'h20;
DFS[16'h0D88] = 8'h95;
DFS[16'h0D89] = 8'h06;
DFS[16'h0D8A] = 8'hBD;
DFS[16'h0D8B] = 8'h00;
DFS[16'h0D8C] = 8'h07;
DFS[16'h0D8D] = 8'h20;
DFS[16'h0D8E] = 8'h95;
DFS[16'h0D8F] = 8'h06;
DFS[16'h0D90] = 8'hE8;
DFS[16'h0D91] = 8'hC9;
DFS[16'h0D92] = 8'h0D;
DFS[16'h0D93] = 8'hD0;
DFS[16'h0D94] = 8'hF5;
DFS[16'h0D95] = 8'h4C;
DFS[16'h0D96] = 8'h36;
DFS[16'h0D97] = 8'h00;
DFS[16'h0D98] = 8'h2C;
DFS[16'h0D99] = 8'hE2;
DFS[16'h0D9A] = 8'hFE;
DFS[16'h0D9B] = 8'h50;
DFS[16'h0D9C] = 8'hFB;
DFS[16'h0D9D] = 8'h8D;
DFS[16'h0D9E] = 8'hE3;
DFS[16'h0D9F] = 8'hFE;
DFS[16'h0DA0] = 8'h60;
DFS[16'h0DA1] = 8'h2C;
DFS[16'h0DA2] = 8'hE6;
DFS[16'h0DA3] = 8'hFE;
DFS[16'h0DA4] = 8'h50;
DFS[16'h0DA5] = 8'hFB;
DFS[16'h0DA6] = 8'h8D;
DFS[16'h0DA7] = 8'hE7;
DFS[16'h0DA8] = 8'hFE;
DFS[16'h0DA9] = 8'h60;
DFS[16'h0DAA] = 8'hA5;
DFS[16'h0DAB] = 8'hFF;
DFS[16'h0DAC] = 8'h38;
DFS[16'h0DAD] = 8'h6A;
DFS[16'h0DAE] = 8'h30;
DFS[16'h0DAF] = 8'h0F;
DFS[16'h0DB0] = 8'h48;
DFS[16'h0DB1] = 8'hA9;
DFS[16'h0DB2] = 8'h00;
DFS[16'h0DB3] = 8'h20;
DFS[16'h0DB4] = 8'hBC;
DFS[16'h0DB5] = 8'h06;
DFS[16'h0DB6] = 8'h98;
DFS[16'h0DB7] = 8'h20;
DFS[16'h0DB8] = 8'hBC;
DFS[16'h0DB9] = 8'h06;
DFS[16'h0DBA] = 8'h8A;
DFS[16'h0DBB] = 8'h20;
DFS[16'h0DBC] = 8'hBC;
DFS[16'h0DBD] = 8'h06;
DFS[16'h0DBE] = 8'h68;
DFS[16'h0DBF] = 8'h2C;
DFS[16'h0DC0] = 8'hE0;
DFS[16'h0DC1] = 8'hFE;
DFS[16'h0DC2] = 8'h50;
DFS[16'h0DC3] = 8'hFB;
DFS[16'h0DC4] = 8'h8D;
DFS[16'h0DC5] = 8'hE1;
DFS[16'h0DC6] = 8'hFE;
DFS[16'h0DC7] = 8'h60;
DFS[16'h0DC8] = 8'h2C;
DFS[16'h0DC9] = 8'hE2;
DFS[16'h0DCA] = 8'hFE;
DFS[16'h0DCB] = 8'h10;
DFS[16'h0DCC] = 8'hFB;
DFS[16'h0DCD] = 8'hAD;
DFS[16'h0DCE] = 8'hE3;
DFS[16'h0DCF] = 8'hFE;
DFS[16'h0DD0] = 8'h60;
DFS[16'h0DD1] = 8'h00;
DFS[16'h0DD2] = 8'h00;
DFS[16'h0DD3] = 8'h00;
DFS[16'h0DD4] = 8'h00;
DFS[16'h0DD5] = 8'h00;
DFS[16'h0DD6] = 8'h00;
DFS[16'h0DD7] = 8'h00;
DFS[16'h0DD8] = 8'h00;
DFS[16'h0DD9] = 8'h00;
DFS[16'h0DDA] = 8'h00;
DFS[16'h0DDB] = 8'h00;
DFS[16'h0DDC] = 8'h00;
DFS[16'h0DDD] = 8'hA2;
DFS[16'h0DDE] = 8'h11;
DFS[16'h0DDF] = 8'hA0;
DFS[16'h0DE0] = 8'h15;
DFS[16'h0DE1] = 8'h60;
DFS[16'h0DE2] = 8'h20;
DFS[16'h0DE3] = 8'hE1;
DFS[16'h0DE4] = 8'h83;
DFS[16'h0DE5] = 8'hA9;
DFS[16'h0DE6] = 8'h77;
DFS[16'h0DE7] = 8'h4C;
DFS[16'h0DE8] = 8'hF4;
DFS[16'h0DE9] = 8'hFF;
DFS[16'h0DEA] = 8'h20;
DFS[16'h0DEB] = 8'hE2;
DFS[16'h0DEC] = 8'h8D;
DFS[16'h0DED] = 8'hA9;
DFS[16'h0DEE] = 8'h00;
DFS[16'h0DEF] = 8'h18;
DFS[16'h0DF0] = 8'h69;
DFS[16'h0DF1] = 8'h20;
DFS[16'h0DF2] = 8'hF0;
DFS[16'h0DF3] = 8'hED;
DFS[16'h0DF4] = 8'hA8;
DFS[16'h0DF5] = 8'h20;
DFS[16'h0DF6] = 8'h05;
DFS[16'h0DF7] = 8'h8E;
DFS[16'h0DF8] = 8'hD0;
DFS[16'h0DF9] = 8'hF5;
DFS[16'h0DFA] = 8'h98;
DFS[16'h0DFB] = 8'hF0;
DFS[16'h0DFC] = 8'hED;
DFS[16'h0DFD] = 8'h20;
DFS[16'h0DFE] = 8'h7B;
DFS[16'h0DFF] = 8'h90;
DFS[16'h0E00] = 8'h90;
DFS[16'h0E01] = 8'h03;
DFS[16'h0E02] = 8'h4C;
DFS[16'h0E03] = 8'hAD;
DFS[16'h0E04] = 8'h90;
DFS[16'h0E05] = 8'h48;
DFS[16'h0E06] = 8'h20;
DFS[16'h0E07] = 8'h51;
DFS[16'h0E08] = 8'h90;
DFS[16'h0E09] = 8'hB0;
DFS[16'h0E0A] = 8'h45;
DFS[16'h0E0B] = 8'hB9;
DFS[16'h0E0C] = 8'h1B;
DFS[16'h0E0D] = 8'h11;
DFS[16'h0E0E] = 8'h49;
DFS[16'h0E0F] = 8'hFF;
DFS[16'h0E10] = 8'h2D;
DFS[16'h0E11] = 8'hC0;
DFS[16'h0E12] = 8'h10;
DFS[16'h0E13] = 8'h8D;
DFS[16'h0E14] = 8'hC0;
DFS[16'h0E15] = 8'h10;
DFS[16'h0E16] = 8'hB9;
DFS[16'h0E17] = 8'h17;
DFS[16'h0E18] = 8'h11;
DFS[16'h0E19] = 8'h29;
DFS[16'h0E1A] = 8'h60;
DFS[16'h0E1B] = 8'hF0;
DFS[16'h0E1C] = 8'h33;
DFS[16'h0E1D] = 8'h20;
DFS[16'h0E1E] = 8'h55;
DFS[16'h0E1F] = 8'h8E;
DFS[16'h0E20] = 8'hB9;
DFS[16'h0E21] = 8'h17;
DFS[16'h0E22] = 8'h11;
DFS[16'h0E23] = 8'h29;
DFS[16'h0E24] = 8'h20;
DFS[16'h0E25] = 8'hF0;
DFS[16'h0E26] = 8'h26;
DFS[16'h0E27] = 8'hAE;
DFS[16'h0E28] = 8'hC4;
DFS[16'h0E29] = 8'h10;
DFS[16'h0E2A] = 8'hB9;
DFS[16'h0E2B] = 8'h14;
DFS[16'h0E2C] = 8'h11;
DFS[16'h0E2D] = 8'h9D;
DFS[16'h0E2E] = 8'h0C;
DFS[16'h0E2F] = 8'h0F;
DFS[16'h0E30] = 8'hB9;
DFS[16'h0E31] = 8'h15;
DFS[16'h0E32] = 8'h11;
DFS[16'h0E33] = 8'h9D;
DFS[16'h0E34] = 8'h0D;
DFS[16'h0E35] = 8'h0F;
DFS[16'h0E36] = 8'hB9;
DFS[16'h0E37] = 8'h16;
DFS[16'h0E38] = 8'h11;
DFS[16'h0E39] = 8'h20;
DFS[16'h0E3A] = 8'h0B;
DFS[16'h0E3B] = 8'h82;
DFS[16'h0E3C] = 8'h5D;
DFS[16'h0E3D] = 8'h0E;
DFS[16'h0E3E] = 8'h0F;
DFS[16'h0E3F] = 8'h29;
DFS[16'h0E40] = 8'h30;
DFS[16'h0E41] = 8'h5D;
DFS[16'h0E42] = 8'h0E;
DFS[16'h0E43] = 8'h0F;
DFS[16'h0E44] = 8'h9D;
DFS[16'h0E45] = 8'h0E;
DFS[16'h0E46] = 8'h0F;
DFS[16'h0E47] = 8'h20;
DFS[16'h0E48] = 8'hB4;
DFS[16'h0E49] = 8'h8A;
DFS[16'h0E4A] = 8'hAC;
DFS[16'h0E4B] = 8'hC2;
DFS[16'h0E4C] = 8'h10;
DFS[16'h0E4D] = 8'h20;
DFS[16'h0E4E] = 8'h4B;
DFS[16'h0E4F] = 8'h91;
DFS[16'h0E50] = 8'hAE;
DFS[16'h0E51] = 8'hC6;
DFS[16'h0E52] = 8'h10;
DFS[16'h0E53] = 8'h68;
DFS[16'h0E54] = 8'h60;
DFS[16'h0E55] = 8'h20;
DFS[16'h0E56] = 8'h83;
DFS[16'h0E57] = 8'h8E;
DFS[16'h0E58] = 8'hA2;
DFS[16'h0E59] = 8'h07;
DFS[16'h0E5A] = 8'hB9;
DFS[16'h0E5B] = 8'h0C;
DFS[16'h0E5C] = 8'h11;
DFS[16'h0E5D] = 8'h95;
DFS[16'h0E5E] = 8'hC6;
DFS[16'h0E5F] = 8'h88;
DFS[16'h0E60] = 8'h88;
DFS[16'h0E61] = 8'hCA;
DFS[16'h0E62] = 8'hD0;
DFS[16'h0E63] = 8'hF6;
DFS[16'h0E64] = 8'h20;
DFS[16'h0E65] = 8'h96;
DFS[16'h0E66] = 8'h82;
DFS[16'h0E67] = 8'h90;
DFS[16'h0E68] = 8'h27;
DFS[16'h0E69] = 8'h8C;
DFS[16'h0E6A] = 8'hC4;
DFS[16'h0E6B] = 8'h10;
DFS[16'h0E6C] = 8'hB9;
DFS[16'h0E6D] = 8'h0E;
DFS[16'h0E6E] = 8'h0F;
DFS[16'h0E6F] = 8'hBE;
DFS[16'h0E70] = 8'h0F;
DFS[16'h0E71] = 8'h0F;
DFS[16'h0E72] = 8'hAC;
DFS[16'h0E73] = 8'hC2;
DFS[16'h0E74] = 8'h10;
DFS[16'h0E75] = 8'h59;
DFS[16'h0E76] = 8'h0D;
DFS[16'h0E77] = 8'h11;
DFS[16'h0E78] = 8'h29;
DFS[16'h0E79] = 8'h03;
DFS[16'h0E7A] = 8'hD0;
DFS[16'h0E7B] = 8'h14;
DFS[16'h0E7C] = 8'h8A;
DFS[16'h0E7D] = 8'hD9;
DFS[16'h0E7E] = 8'h0F;
DFS[16'h0E7F] = 8'h11;
DFS[16'h0E80] = 8'hD0;
DFS[16'h0E81] = 8'h0E;
DFS[16'h0E82] = 8'h60;
DFS[16'h0E83] = 8'hB9;
DFS[16'h0E84] = 8'h0E;
DFS[16'h0E85] = 8'h11;
DFS[16'h0E86] = 8'h29;
DFS[16'h0E87] = 8'h7F;
DFS[16'h0E88] = 8'h85;
DFS[16'h0E89] = 8'hCE;
DFS[16'h0E8A] = 8'hB9;
DFS[16'h0E8B] = 8'h17;
DFS[16'h0E8C] = 8'h11;
DFS[16'h0E8D] = 8'h4C;
DFS[16'h0E8E] = 8'h7E;
DFS[16'h0E8F] = 8'h87;
DFS[16'h0E90] = 8'h4C;
DFS[16'h0E91] = 8'hAF;
DFS[16'h0E92] = 8'h81;
DFS[16'h0E93] = 8'hC9;
DFS[16'h0E94] = 8'h00;
DFS[16'h0E95] = 8'hD0;
DFS[16'h0E96] = 8'h06;
DFS[16'h0E97] = 8'h20;
DFS[16'h0E98] = 8'hE1;
DFS[16'h0E99] = 8'h83;
DFS[16'h0E9A] = 8'h4C;
DFS[16'h0E9B] = 8'hFA;
DFS[16'h0E9C] = 8'h8D;
DFS[16'h0E9D] = 8'h20;
DFS[16'h0E9E] = 8'h11;
DFS[16'h0E9F] = 8'h84;
DFS[16'h0EA0] = 8'h86;
DFS[16'h0EA1] = 8'hBC;
DFS[16'h0EA2] = 8'h84;
DFS[16'h0EA3] = 8'hBD;
DFS[16'h0EA4] = 8'h85;
DFS[16'h0EA5] = 8'hB4;
DFS[16'h0EA6] = 8'h24;
DFS[16'h0EA7] = 8'hB4;
DFS[16'h0EA8] = 8'h08;
DFS[16'h0EA9] = 8'h20;
DFS[16'h0EAA] = 8'h06;
DFS[16'h0EAB] = 8'h81;
DFS[16'h0EAC] = 8'h20;
DFS[16'h0EAD] = 8'h96;
DFS[16'h0EAE] = 8'h82;
DFS[16'h0EAF] = 8'hB0;
DFS[16'h0EB0] = 8'h1A;
DFS[16'h0EB1] = 8'h28;
DFS[16'h0EB2] = 8'h50;
DFS[16'h0EB3] = 8'h03;
DFS[16'h0EB4] = 8'hA9;
DFS[16'h0EB5] = 8'h00;
DFS[16'h0EB6] = 8'h60;
DFS[16'h0EB7] = 8'h08;
DFS[16'h0EB8] = 8'hA9;
DFS[16'h0EB9] = 8'h00;
DFS[16'h0EBA] = 8'hA2;
DFS[16'h0EBB] = 8'h07;
DFS[16'h0EBC] = 8'h95;
DFS[16'h0EBD] = 8'hBE;
DFS[16'h0EBE] = 8'h9D;
DFS[16'h0EBF] = 8'h74;
DFS[16'h0EC0] = 8'h10;
DFS[16'h0EC1] = 8'hCA;
DFS[16'h0EC2] = 8'h10;
DFS[16'h0EC3] = 8'hF8;
DFS[16'h0EC4] = 8'hA9;
DFS[16'h0EC5] = 8'h40;
DFS[16'h0EC6] = 8'h85;
DFS[16'h0EC7] = 8'hC5;
DFS[16'h0EC8] = 8'h20;
DFS[16'h0EC9] = 8'h61;
DFS[16'h0ECA] = 8'h89;
DFS[16'h0ECB] = 8'h28;
DFS[16'h0ECC] = 8'h08;
DFS[16'h0ECD] = 8'h70;
DFS[16'h0ECE] = 8'h03;
DFS[16'h0ECF] = 8'h20;
DFS[16'h0ED0] = 8'h3C;
DFS[16'h0ED1] = 8'h98;
DFS[16'h0ED2] = 8'h20;
DFS[16'h0ED3] = 8'h9E;
DFS[16'h0ED4] = 8'h8F;
DFS[16'h0ED5] = 8'h90;
DFS[16'h0ED6] = 8'h0E;
DFS[16'h0ED7] = 8'hB9;
DFS[16'h0ED8] = 8'h0C;
DFS[16'h0ED9] = 8'h11;
DFS[16'h0EDA] = 8'h10;
DFS[16'h0EDB] = 8'h26;
DFS[16'h0EDC] = 8'h24;
DFS[16'h0EDD] = 8'hB4;
DFS[16'h0EDE] = 8'h30;
DFS[16'h0EDF] = 8'h22;
DFS[16'h0EE0] = 8'h20;
DFS[16'h0EE1] = 8'h99;
DFS[16'h0EE2] = 8'h8F;
DFS[16'h0EE3] = 8'hB0;
DFS[16'h0EE4] = 8'hF2;
DFS[16'h0EE5] = 8'hAC;
DFS[16'h0EE6] = 8'hC2;
DFS[16'h0EE7] = 8'h10;
DFS[16'h0EE8] = 8'hD0;
DFS[16'h0EE9] = 8'h21;
DFS[16'h0EEA] = 8'h20;
DFS[16'h0EEB] = 8'h33;
DFS[16'h0EEC] = 8'h80;
DFS[16'h0EED] = 8'hC0;
DFS[16'h0EEE] = 8'h54;
DFS[16'h0EEF] = 8'h6F;
DFS[16'h0EF0] = 8'h6F;
DFS[16'h0EF1] = 8'h20;
DFS[16'h0EF2] = 8'h6D;
DFS[16'h0EF3] = 8'h61;
DFS[16'h0EF4] = 8'h6E;
DFS[16'h0EF5] = 8'h79;
DFS[16'h0EF6] = 8'h20;
DFS[16'h0EF7] = 8'h66;
DFS[16'h0EF8] = 8'h69;
DFS[16'h0EF9] = 8'h6C;
DFS[16'h0EFA] = 8'h65;
DFS[16'h0EFB] = 8'h73;
DFS[16'h0EFC] = 8'h20;
DFS[16'h0EFD] = 8'h6F;
DFS[16'h0EFE] = 8'h70;
DFS[16'h0EFF] = 8'h65;
DFS[16'h0F00] = 8'h6E;
DFS[16'h0F01] = 8'h00;
DFS[16'h0F02] = 8'h20;
DFS[16'h0F03] = 8'h2B;
DFS[16'h0F04] = 8'h80;
DFS[16'h0F05] = 8'hC2;
DFS[16'h0F06] = 8'h6F;
DFS[16'h0F07] = 8'h70;
DFS[16'h0F08] = 8'h65;
DFS[16'h0F09] = 8'h6E;
DFS[16'h0F0A] = 8'h00;
DFS[16'h0F0B] = 8'hA9;
DFS[16'h0F0C] = 8'h08;
DFS[16'h0F0D] = 8'h8D;
DFS[16'h0F0E] = 8'hC5;
DFS[16'h0F0F] = 8'h10;
DFS[16'h0F10] = 8'hBD;
DFS[16'h0F11] = 8'h08;
DFS[16'h0F12] = 8'h0E;
DFS[16'h0F13] = 8'h99;
DFS[16'h0F14] = 8'h00;
DFS[16'h0F15] = 8'h11;
DFS[16'h0F16] = 8'hC8;
DFS[16'h0F17] = 8'hBD;
DFS[16'h0F18] = 8'h08;
DFS[16'h0F19] = 8'h0F;
DFS[16'h0F1A] = 8'h99;
DFS[16'h0F1B] = 8'h00;
DFS[16'h0F1C] = 8'h11;
DFS[16'h0F1D] = 8'hC8;
DFS[16'h0F1E] = 8'hE8;
DFS[16'h0F1F] = 8'hCE;
DFS[16'h0F20] = 8'hC5;
DFS[16'h0F21] = 8'h10;
DFS[16'h0F22] = 8'hD0;
DFS[16'h0F23] = 8'hEC;
DFS[16'h0F24] = 8'hA2;
DFS[16'h0F25] = 8'h10;
DFS[16'h0F26] = 8'hA9;
DFS[16'h0F27] = 8'h00;
DFS[16'h0F28] = 8'h99;
DFS[16'h0F29] = 8'h00;
DFS[16'h0F2A] = 8'h11;
DFS[16'h0F2B] = 8'hC8;
DFS[16'h0F2C] = 8'hCA;
DFS[16'h0F2D] = 8'hD0;
DFS[16'h0F2E] = 8'hF9;
DFS[16'h0F2F] = 8'hAD;
DFS[16'h0F30] = 8'hC2;
DFS[16'h0F31] = 8'h10;
DFS[16'h0F32] = 8'hA8;
DFS[16'h0F33] = 8'h20;
DFS[16'h0F34] = 8'h04;
DFS[16'h0F35] = 8'h82;
DFS[16'h0F36] = 8'h69;
DFS[16'h0F37] = 8'h11;
DFS[16'h0F38] = 8'h99;
DFS[16'h0F39] = 8'h13;
DFS[16'h0F3A] = 8'h11;
DFS[16'h0F3B] = 8'hAD;
DFS[16'h0F3C] = 8'hC1;
DFS[16'h0F3D] = 8'h10;
DFS[16'h0F3E] = 8'h99;
DFS[16'h0F3F] = 8'h1B;
DFS[16'h0F40] = 8'h11;
DFS[16'h0F41] = 8'h0D;
DFS[16'h0F42] = 8'hC0;
DFS[16'h0F43] = 8'h10;
DFS[16'h0F44] = 8'h8D;
DFS[16'h0F45] = 8'hC0;
DFS[16'h0F46] = 8'h10;
DFS[16'h0F47] = 8'hB9;
DFS[16'h0F48] = 8'h09;
DFS[16'h0F49] = 8'h11;
DFS[16'h0F4A] = 8'h69;
DFS[16'h0F4B] = 8'hFF;
DFS[16'h0F4C] = 8'hB9;
DFS[16'h0F4D] = 8'h0B;
DFS[16'h0F4E] = 8'h11;
DFS[16'h0F4F] = 8'h69;
DFS[16'h0F50] = 8'h00;
DFS[16'h0F51] = 8'h99;
DFS[16'h0F52] = 8'h19;
DFS[16'h0F53] = 8'h11;
DFS[16'h0F54] = 8'hB9;
DFS[16'h0F55] = 8'h0D;
DFS[16'h0F56] = 8'h11;
DFS[16'h0F57] = 8'h09;
DFS[16'h0F58] = 8'h0F;
DFS[16'h0F59] = 8'h69;
DFS[16'h0F5A] = 8'h00;
DFS[16'h0F5B] = 8'h20;
DFS[16'h0F5C] = 8'hFD;
DFS[16'h0F5D] = 8'h81;
DFS[16'h0F5E] = 8'h99;
DFS[16'h0F5F] = 8'h1A;
DFS[16'h0F60] = 8'h11;
DFS[16'h0F61] = 8'h28;
DFS[16'h0F62] = 8'h50;
DFS[16'h0F63] = 8'h2E;
DFS[16'h0F64] = 8'h30;
DFS[16'h0F65] = 8'h08;
DFS[16'h0F66] = 8'hA9;
DFS[16'h0F67] = 8'h80;
DFS[16'h0F68] = 8'h19;
DFS[16'h0F69] = 8'h0C;
DFS[16'h0F6A] = 8'h11;
DFS[16'h0F6B] = 8'h99;
DFS[16'h0F6C] = 8'h0C;
DFS[16'h0F6D] = 8'h11;
DFS[16'h0F6E] = 8'hB9;
DFS[16'h0F6F] = 8'h09;
DFS[16'h0F70] = 8'h11;
DFS[16'h0F71] = 8'h99;
DFS[16'h0F72] = 8'h14;
DFS[16'h0F73] = 8'h11;
DFS[16'h0F74] = 8'hB9;
DFS[16'h0F75] = 8'h0B;
DFS[16'h0F76] = 8'h11;
DFS[16'h0F77] = 8'h99;
DFS[16'h0F78] = 8'h15;
DFS[16'h0F79] = 8'h11;
DFS[16'h0F7A] = 8'hB9;
DFS[16'h0F7B] = 8'h0D;
DFS[16'h0F7C] = 8'h11;
DFS[16'h0F7D] = 8'h20;
DFS[16'h0F7E] = 8'hFD;
DFS[16'h0F7F] = 8'h81;
DFS[16'h0F80] = 8'h99;
DFS[16'h0F81] = 8'h16;
DFS[16'h0F82] = 8'h11;
DFS[16'h0F83] = 8'hA5;
DFS[16'h0F84] = 8'hCF;
DFS[16'h0F85] = 8'h19;
DFS[16'h0F86] = 8'h17;
DFS[16'h0F87] = 8'h11;
DFS[16'h0F88] = 8'h99;
DFS[16'h0F89] = 8'h17;
DFS[16'h0F8A] = 8'h11;
DFS[16'h0F8B] = 8'h98;
DFS[16'h0F8C] = 8'h20;
DFS[16'h0F8D] = 8'h04;
DFS[16'h0F8E] = 8'h82;
DFS[16'h0F8F] = 8'h09;
DFS[16'h0F90] = 8'h10;
DFS[16'h0F91] = 8'h60;
DFS[16'h0F92] = 8'hA9;
DFS[16'h0F93] = 8'h20;
DFS[16'h0F94] = 8'h99;
DFS[16'h0F95] = 8'h17;
DFS[16'h0F96] = 8'h11;
DFS[16'h0F97] = 8'hD0;
DFS[16'h0F98] = 8'hEA;
DFS[16'h0F99] = 8'h8A;
DFS[16'h0F9A] = 8'h48;
DFS[16'h0F9B] = 8'h4C;
DFS[16'h0F9C] = 8'hDD;
DFS[16'h0F9D] = 8'h8F;
DFS[16'h0F9E] = 8'hA9;
DFS[16'h0F9F] = 8'h00;
DFS[16'h0FA0] = 8'h8D;
DFS[16'h0FA1] = 8'hC2;
DFS[16'h0FA2] = 8'h10;
DFS[16'h0FA3] = 8'hA9;
DFS[16'h0FA4] = 8'h08;
DFS[16'h0FA5] = 8'h85;
DFS[16'h0FA6] = 8'hB5;
DFS[16'h0FA7] = 8'h98;
DFS[16'h0FA8] = 8'hAA;
DFS[16'h0FA9] = 8'hA0;
DFS[16'h0FAA] = 8'hA0;
DFS[16'h0FAB] = 8'h84;
DFS[16'h0FAC] = 8'hB3;
DFS[16'h0FAD] = 8'h8A;
DFS[16'h0FAE] = 8'h48;
DFS[16'h0FAF] = 8'hA9;
DFS[16'h0FB0] = 8'h08;
DFS[16'h0FB1] = 8'h85;
DFS[16'h0FB2] = 8'hB2;
DFS[16'h0FB3] = 8'hA5;
DFS[16'h0FB4] = 8'hB5;
DFS[16'h0FB5] = 8'h2C;
DFS[16'h0FB6] = 8'hC0;
DFS[16'h0FB7] = 8'h10;
DFS[16'h0FB8] = 8'hF0;
DFS[16'h0FB9] = 8'h1D;
DFS[16'h0FBA] = 8'hB9;
DFS[16'h0FBB] = 8'h17;
DFS[16'h0FBC] = 8'h11;
DFS[16'h0FBD] = 8'h45;
DFS[16'h0FBE] = 8'hCF;
DFS[16'h0FBF] = 8'h29;
DFS[16'h0FC0] = 8'h03;
DFS[16'h0FC1] = 8'hD0;
DFS[16'h0FC2] = 8'h1A;
DFS[16'h0FC3] = 8'hBD;
DFS[16'h0FC4] = 8'h08;
DFS[16'h0FC5] = 8'h0E;
DFS[16'h0FC6] = 8'h59;
DFS[16'h0FC7] = 8'h00;
DFS[16'h0FC8] = 8'h11;
DFS[16'h0FC9] = 8'h29;
DFS[16'h0FCA] = 8'h7F;
DFS[16'h0FCB] = 8'hD0;
DFS[16'h0FCC] = 8'h10;
DFS[16'h0FCD] = 8'hE8;
DFS[16'h0FCE] = 8'hC8;
DFS[16'h0FCF] = 8'hC8;
DFS[16'h0FD0] = 8'hC6;
DFS[16'h0FD1] = 8'hB2;
DFS[16'h0FD2] = 8'hD0;
DFS[16'h0FD3] = 8'hEF;
DFS[16'h0FD4] = 8'h38;
DFS[16'h0FD5] = 8'hB0;
DFS[16'h0FD6] = 8'h10;
DFS[16'h0FD7] = 8'h8C;
DFS[16'h0FD8] = 8'hC2;
DFS[16'h0FD9] = 8'h10;
DFS[16'h0FDA] = 8'h8D;
DFS[16'h0FDB] = 8'hC1;
DFS[16'h0FDC] = 8'h10;
DFS[16'h0FDD] = 8'h38;
DFS[16'h0FDE] = 8'hA5;
DFS[16'h0FDF] = 8'hB3;
DFS[16'h0FE0] = 8'hE9;
DFS[16'h0FE1] = 8'h20;
DFS[16'h0FE2] = 8'h85;
DFS[16'h0FE3] = 8'hB3;
DFS[16'h0FE4] = 8'h06;
DFS[16'h0FE5] = 8'hB5;
DFS[16'h0FE6] = 8'h18;
DFS[16'h0FE7] = 8'h68;
DFS[16'h0FE8] = 8'hAA;
DFS[16'h0FE9] = 8'hA4;
DFS[16'h0FEA] = 8'hB3;
DFS[16'h0FEB] = 8'hA5;
DFS[16'h0FEC] = 8'hB5;
DFS[16'h0FED] = 8'hB0;
DFS[16'h0FEE] = 8'h02;
DFS[16'h0FEF] = 8'hD0;
DFS[16'h0FF0] = 8'hBA;
DFS[16'h0FF1] = 8'h60;
DFS[16'h0FF2] = 8'hAD;
DFS[16'h0FF3] = 8'hC0;
DFS[16'h0FF4] = 8'h10;
DFS[16'h0FF5] = 8'h48;
DFS[16'h0FF6] = 8'h20;
DFS[16'h0FF7] = 8'hED;
DFS[16'h0FF8] = 8'h8D;
DFS[16'h0FF9] = 8'hF0;
DFS[16'h0FFA] = 8'h07;
DFS[16'h0FFB] = 8'hAD;
DFS[16'h0FFC] = 8'hC0;
DFS[16'h0FFD] = 8'h10;
DFS[16'h0FFE] = 8'h48;
DFS[16'h0FFF] = 8'h20;
DFS[16'h1000] = 8'hFA;
DFS[16'h1001] = 8'h8D;
DFS[16'h1002] = 8'h68;
DFS[16'h1003] = 8'h8D;
DFS[16'h1004] = 8'hC0;
DFS[16'h1005] = 8'h10;
DFS[16'h1006] = 8'h60;
DFS[16'h1007] = 8'hC0;
DFS[16'h1008] = 8'h00;
DFS[16'h1009] = 8'hF0;
DFS[16'h100A] = 8'h11;
DFS[16'h100B] = 8'h20;
DFS[16'h100C] = 8'hE1;
DFS[16'h100D] = 8'h83;
DFS[16'h100E] = 8'hC9;
DFS[16'h100F] = 8'hFF;
DFS[16'h1010] = 8'hF0;
DFS[16'h1011] = 8'hE9;
DFS[16'h1012] = 8'hC9;
DFS[16'h1013] = 8'h03;
DFS[16'h1014] = 8'hB0;
DFS[16'h1015] = 8'h17;
DFS[16'h1016] = 8'h4A;
DFS[16'h1017] = 8'h90;
DFS[16'h1018] = 8'h15;
DFS[16'h1019] = 8'h4C;
DFS[16'h101A] = 8'hA7;
DFS[16'h101B] = 8'h92;
DFS[16'h101C] = 8'h20;
DFS[16'h101D] = 8'h11;
DFS[16'h101E] = 8'h84;
DFS[16'h101F] = 8'hA8;
DFS[16'h1020] = 8'hC8;
DFS[16'h1021] = 8'hC0;
DFS[16'h1022] = 8'h03;
DFS[16'h1023] = 8'hB0;
DFS[16'h1024] = 8'h08;
DFS[16'h1025] = 8'hB9;
DFS[16'h1026] = 8'h81;
DFS[16'h1027] = 8'h99;
DFS[16'h1028] = 8'h48;
DFS[16'h1029] = 8'hB9;
DFS[16'h102A] = 8'h7E;
DFS[16'h102B] = 8'h99;
DFS[16'h102C] = 8'h48;
DFS[16'h102D] = 8'h60;
DFS[16'h102E] = 8'h20;
DFS[16'h102F] = 8'hE1;
DFS[16'h1030] = 8'h83;
DFS[16'h1031] = 8'h20;
DFS[16'h1032] = 8'hA5;
DFS[16'h1033] = 8'h90;
DFS[16'h1034] = 8'h8C;
DFS[16'h1035] = 8'hC2;
DFS[16'h1036] = 8'h10;
DFS[16'h1037] = 8'h0A;
DFS[16'h1038] = 8'h0A;
DFS[16'h1039] = 8'h6D;
DFS[16'h103A] = 8'hC2;
DFS[16'h103B] = 8'h10;
DFS[16'h103C] = 8'hA8;
DFS[16'h103D] = 8'hB9;
DFS[16'h103E] = 8'h10;
DFS[16'h103F] = 8'h11;
DFS[16'h1040] = 8'h95;
DFS[16'h1041] = 8'h00;
DFS[16'h1042] = 8'hB9;
DFS[16'h1043] = 8'h11;
DFS[16'h1044] = 8'h11;
DFS[16'h1045] = 8'h95;
DFS[16'h1046] = 8'h01;
DFS[16'h1047] = 8'hB9;
DFS[16'h1048] = 8'h12;
DFS[16'h1049] = 8'h11;
DFS[16'h104A] = 8'h95;
DFS[16'h104B] = 8'h02;
DFS[16'h104C] = 8'hA9;
DFS[16'h104D] = 8'h00;
DFS[16'h104E] = 8'h95;
DFS[16'h104F] = 8'h03;
DFS[16'h1050] = 8'h60;
DFS[16'h1051] = 8'h48;
DFS[16'h1052] = 8'h8E;
DFS[16'h1053] = 8'hC6;
DFS[16'h1054] = 8'h10;
DFS[16'h1055] = 8'h98;
DFS[16'h1056] = 8'h29;
DFS[16'h1057] = 8'hE0;
DFS[16'h1058] = 8'h8D;
DFS[16'h1059] = 8'hC2;
DFS[16'h105A] = 8'h10;
DFS[16'h105B] = 8'hF0;
DFS[16'h105C] = 8'h13;
DFS[16'h105D] = 8'h20;
DFS[16'h105E] = 8'h04;
DFS[16'h105F] = 8'h82;
DFS[16'h1060] = 8'hA8;
DFS[16'h1061] = 8'hA9;
DFS[16'h1062] = 8'h00;
DFS[16'h1063] = 8'h38;
DFS[16'h1064] = 8'h6A;
DFS[16'h1065] = 8'h88;
DFS[16'h1066] = 8'hD0;
DFS[16'h1067] = 8'hFC;
DFS[16'h1068] = 8'hAC;
DFS[16'h1069] = 8'hC2;
DFS[16'h106A] = 8'h10;
DFS[16'h106B] = 8'h2C;
DFS[16'h106C] = 8'hC0;
DFS[16'h106D] = 8'h10;
DFS[16'h106E] = 8'hD0;
DFS[16'h106F] = 8'h03;
DFS[16'h1070] = 8'h68;
DFS[16'h1071] = 8'h38;
DFS[16'h1072] = 8'h60;
DFS[16'h1073] = 8'h68;
DFS[16'h1074] = 8'h18;
DFS[16'h1075] = 8'h60;
DFS[16'h1076] = 8'h48;
DFS[16'h1077] = 8'h8A;
DFS[16'h1078] = 8'h4C;
DFS[16'h1079] = 8'h7D;
DFS[16'h107A] = 8'h90;
DFS[16'h107B] = 8'h48;
DFS[16'h107C] = 8'h98;
DFS[16'h107D] = 8'hC9;
DFS[16'h107E] = 8'h10;
DFS[16'h107F] = 8'h90;
DFS[16'h1080] = 8'h04;
DFS[16'h1081] = 8'hC9;
DFS[16'h1082] = 8'h18;
DFS[16'h1083] = 8'h90;
DFS[16'h1084] = 8'h02;
DFS[16'h1085] = 8'hA9;
DFS[16'h1086] = 8'h08;
DFS[16'h1087] = 8'h20;
DFS[16'h1088] = 8'h0A;
DFS[16'h1089] = 8'h82;
DFS[16'h108A] = 8'hA8;
DFS[16'h108B] = 8'h68;
DFS[16'h108C] = 8'h60;
DFS[16'h108D] = 8'h48;
DFS[16'h108E] = 8'h98;
DFS[16'h108F] = 8'h48;
DFS[16'h1090] = 8'h8A;
DFS[16'h1091] = 8'hA8;
DFS[16'h1092] = 8'h20;
DFS[16'h1093] = 8'hA5;
DFS[16'h1094] = 8'h90;
DFS[16'h1095] = 8'h98;
DFS[16'h1096] = 8'h20;
DFS[16'h1097] = 8'hF8;
DFS[16'h1098] = 8'h92;
DFS[16'h1099] = 8'hD0;
DFS[16'h109A] = 8'h04;
DFS[16'h109B] = 8'hA2;
DFS[16'h109C] = 8'hFF;
DFS[16'h109D] = 8'hD0;
DFS[16'h109E] = 8'h02;
DFS[16'h109F] = 8'hA2;
DFS[16'h10A0] = 8'h00;
DFS[16'h10A1] = 8'h68;
DFS[16'h10A2] = 8'hA8;
DFS[16'h10A3] = 8'h68;
DFS[16'h10A4] = 8'h60;
DFS[16'h10A5] = 8'h20;
DFS[16'h10A6] = 8'h7B;
DFS[16'h10A7] = 8'h90;
DFS[16'h10A8] = 8'h20;
DFS[16'h10A9] = 8'h51;
DFS[16'h10AA] = 8'h90;
DFS[16'h10AB] = 8'h90;
DFS[16'h10AC] = 8'hF7;
DFS[16'h10AD] = 8'h20;
DFS[16'h10AE] = 8'h33;
DFS[16'h10AF] = 8'h80;
DFS[16'h10B0] = 8'hDE;
DFS[16'h10B1] = 8'h43;
DFS[16'h10B2] = 8'h68;
DFS[16'h10B3] = 8'h61;
DFS[16'h10B4] = 8'h6E;
DFS[16'h10B5] = 8'h6E;
DFS[16'h10B6] = 8'h65;
DFS[16'h10B7] = 8'h6C;
DFS[16'h10B8] = 8'h00;
DFS[16'h10B9] = 8'h20;
DFS[16'h10BA] = 8'h33;
DFS[16'h10BB] = 8'h80;
DFS[16'h10BC] = 8'hDF;
DFS[16'h10BD] = 8'h45;
DFS[16'h10BE] = 8'h4F;
DFS[16'h10BF] = 8'h46;
DFS[16'h10C0] = 8'h00;
DFS[16'h10C1] = 8'h20;
DFS[16'h10C2] = 8'h11;
DFS[16'h10C3] = 8'h84;
DFS[16'h10C4] = 8'h20;
DFS[16'h10C5] = 8'hA5;
DFS[16'h10C6] = 8'h90;
DFS[16'h10C7] = 8'h98;
DFS[16'h10C8] = 8'h20;
DFS[16'h10C9] = 8'hF8;
DFS[16'h10CA] = 8'h92;
DFS[16'h10CB] = 8'hD0;
DFS[16'h10CC] = 8'h13;
DFS[16'h10CD] = 8'hB9;
DFS[16'h10CE] = 8'h17;
DFS[16'h10CF] = 8'h11;
DFS[16'h10D0] = 8'h29;
DFS[16'h10D1] = 8'h10;
DFS[16'h10D2] = 8'hD0;
DFS[16'h10D3] = 8'hE5;
DFS[16'h10D4] = 8'hA9;
DFS[16'h10D5] = 8'h10;
DFS[16'h10D6] = 8'h20;
DFS[16'h10D7] = 8'h3C;
DFS[16'h10D8] = 8'h91;
DFS[16'h10D9] = 8'hAE;
DFS[16'h10DA] = 8'hC6;
DFS[16'h10DB] = 8'h10;
DFS[16'h10DC] = 8'hA9;
DFS[16'h10DD] = 8'hFE;
DFS[16'h10DE] = 8'h38;
DFS[16'h10DF] = 8'h60;
DFS[16'h10E0] = 8'hB9;
DFS[16'h10E1] = 8'h17;
DFS[16'h10E2] = 8'h11;
DFS[16'h10E3] = 8'h30;
DFS[16'h10E4] = 8'h0A;
DFS[16'h10E5] = 8'h20;
DFS[16'h10E6] = 8'h83;
DFS[16'h10E7] = 8'h8E;
DFS[16'h10E8] = 8'h20;
DFS[16'h10E9] = 8'h4B;
DFS[16'h10EA] = 8'h91;
DFS[16'h10EB] = 8'h38;
DFS[16'h10EC] = 8'h20;
DFS[16'h10ED] = 8'h53;
DFS[16'h10EE] = 8'h91;
DFS[16'h10EF] = 8'hB9;
DFS[16'h10F0] = 8'h10;
DFS[16'h10F1] = 8'h11;
DFS[16'h10F2] = 8'h85;
DFS[16'h10F3] = 8'hBC;
DFS[16'h10F4] = 8'hB9;
DFS[16'h10F5] = 8'h13;
DFS[16'h10F6] = 8'h11;
DFS[16'h10F7] = 8'h85;
DFS[16'h10F8] = 8'hBD;
DFS[16'h10F9] = 8'hA0;
DFS[16'h10FA] = 8'h00;
DFS[16'h10FB] = 8'hB1;
DFS[16'h10FC] = 8'hBC;
DFS[16'h10FD] = 8'h48;
DFS[16'h10FE] = 8'hAC;
DFS[16'h10FF] = 8'hC2;
DFS[16'h1100] = 8'h10;
DFS[16'h1101] = 8'hA6;
DFS[16'h1102] = 8'hBC;
DFS[16'h1103] = 8'hE8;
DFS[16'h1104] = 8'h8A;
DFS[16'h1105] = 8'h99;
DFS[16'h1106] = 8'h10;
DFS[16'h1107] = 8'h11;
DFS[16'h1108] = 8'hD0;
DFS[16'h1109] = 8'h14;
DFS[16'h110A] = 8'h18;
DFS[16'h110B] = 8'hB9;
DFS[16'h110C] = 8'h11;
DFS[16'h110D] = 8'h11;
DFS[16'h110E] = 8'h69;
DFS[16'h110F] = 8'h01;
DFS[16'h1110] = 8'h99;
DFS[16'h1111] = 8'h11;
DFS[16'h1112] = 8'h11;
DFS[16'h1113] = 8'hB9;
DFS[16'h1114] = 8'h12;
DFS[16'h1115] = 8'h11;
DFS[16'h1116] = 8'h69;
DFS[16'h1117] = 8'h00;
DFS[16'h1118] = 8'h99;
DFS[16'h1119] = 8'h12;
DFS[16'h111A] = 8'h11;
DFS[16'h111B] = 8'h20;
DFS[16'h111C] = 8'h41;
DFS[16'h111D] = 8'h91;
DFS[16'h111E] = 8'h18;
DFS[16'h111F] = 8'h68;
DFS[16'h1120] = 8'h60;
DFS[16'h1121] = 8'h18;
DFS[16'h1122] = 8'hB9;
DFS[16'h1123] = 8'h0F;
DFS[16'h1124] = 8'h11;
DFS[16'h1125] = 8'h79;
DFS[16'h1126] = 8'h11;
DFS[16'h1127] = 8'h11;
DFS[16'h1128] = 8'h85;
DFS[16'h1129] = 8'hC5;
DFS[16'h112A] = 8'h99;
DFS[16'h112B] = 8'h1C;
DFS[16'h112C] = 8'h11;
DFS[16'h112D] = 8'hB9;
DFS[16'h112E] = 8'h0D;
DFS[16'h112F] = 8'h11;
DFS[16'h1130] = 8'h29;
DFS[16'h1131] = 8'h03;
DFS[16'h1132] = 8'h79;
DFS[16'h1133] = 8'h12;
DFS[16'h1134] = 8'h11;
DFS[16'h1135] = 8'h85;
DFS[16'h1136] = 8'hC4;
DFS[16'h1137] = 8'h99;
DFS[16'h1138] = 8'h1D;
DFS[16'h1139] = 8'h11;
DFS[16'h113A] = 8'hA9;
DFS[16'h113B] = 8'h80;
DFS[16'h113C] = 8'h19;
DFS[16'h113D] = 8'h17;
DFS[16'h113E] = 8'h11;
DFS[16'h113F] = 8'hD0;
DFS[16'h1140] = 8'h05;
DFS[16'h1141] = 8'hA9;
DFS[16'h1142] = 8'h7F;
DFS[16'h1143] = 8'h39;
DFS[16'h1144] = 8'h17;
DFS[16'h1145] = 8'h11;
DFS[16'h1146] = 8'h99;
DFS[16'h1147] = 8'h17;
DFS[16'h1148] = 8'h11;
DFS[16'h1149] = 8'h18;
DFS[16'h114A] = 8'h60;
DFS[16'h114B] = 8'hB9;
DFS[16'h114C] = 8'h17;
DFS[16'h114D] = 8'h11;
DFS[16'h114E] = 8'h29;
DFS[16'h114F] = 8'h40;
DFS[16'h1150] = 8'hF0;
DFS[16'h1151] = 8'h3D;
DFS[16'h1152] = 8'h18;
DFS[16'h1153] = 8'h08;
DFS[16'h1154] = 8'h20;
DFS[16'h1155] = 8'h0B;
DFS[16'h1156] = 8'hB9;
DFS[16'h1157] = 8'hAC;
DFS[16'h1158] = 8'hC2;
DFS[16'h1159] = 8'h10;
DFS[16'h115A] = 8'hB9;
DFS[16'h115B] = 8'h13;
DFS[16'h115C] = 8'h11;
DFS[16'h115D] = 8'h85;
DFS[16'h115E] = 8'hBF;
DFS[16'h115F] = 8'h20;
DFS[16'h1160] = 8'h8D;
DFS[16'h1161] = 8'hA0;
DFS[16'h1162] = 8'hA9;
DFS[16'h1163] = 8'h00;
DFS[16'h1164] = 8'h85;
DFS[16'h1165] = 8'hBE;
DFS[16'h1166] = 8'h85;
DFS[16'h1167] = 8'hC2;
DFS[16'h1168] = 8'hA9;
DFS[16'h1169] = 8'h01;
DFS[16'h116A] = 8'h85;
DFS[16'h116B] = 8'hC3;
DFS[16'h116C] = 8'h28;
DFS[16'h116D] = 8'hB0;
DFS[16'h116E] = 8'h17;
DFS[16'h116F] = 8'hB9;
DFS[16'h1170] = 8'h1C;
DFS[16'h1171] = 8'h11;
DFS[16'h1172] = 8'h85;
DFS[16'h1173] = 8'hC5;
DFS[16'h1174] = 8'hB9;
DFS[16'h1175] = 8'h1D;
DFS[16'h1176] = 8'h11;
DFS[16'h1177] = 8'h85;
DFS[16'h1178] = 8'hC4;
DFS[16'h1179] = 8'h20;
DFS[16'h117A] = 8'h8F;
DFS[16'h117B] = 8'h87;
DFS[16'h117C] = 8'hAC;
DFS[16'h117D] = 8'hC2;
DFS[16'h117E] = 8'h10;
DFS[16'h117F] = 8'hA9;
DFS[16'h1180] = 8'hBF;
DFS[16'h1181] = 8'h20;
DFS[16'h1182] = 8'h43;
DFS[16'h1183] = 8'h91;
DFS[16'h1184] = 8'h90;
DFS[16'h1185] = 8'h06;
DFS[16'h1186] = 8'h20;
DFS[16'h1187] = 8'h21;
DFS[16'h1188] = 8'h91;
DFS[16'h1189] = 8'h20;
DFS[16'h118A] = 8'hC6;
DFS[16'h118B] = 8'h87;
DFS[16'h118C] = 8'hAC;
DFS[16'h118D] = 8'hC2;
DFS[16'h118E] = 8'h10;
DFS[16'h118F] = 8'h60;
DFS[16'h1190] = 8'h4C;
DFS[16'h1191] = 8'hAD;
DFS[16'h1192] = 8'h90;
DFS[16'h1193] = 8'h4C;
DFS[16'h1194] = 8'h41;
DFS[16'h1195] = 8'h98;
DFS[16'h1196] = 8'h20;
DFS[16'h1197] = 8'h2B;
DFS[16'h1198] = 8'h80;
DFS[16'h1199] = 8'hC1;
DFS[16'h119A] = 8'h72;
DFS[16'h119B] = 8'h65;
DFS[16'h119C] = 8'h61;
DFS[16'h119D] = 8'h64;
DFS[16'h119E] = 8'h20;
DFS[16'h119F] = 8'h6F;
DFS[16'h11A0] = 8'h6E;
DFS[16'h11A1] = 8'h6C;
DFS[16'h11A2] = 8'h79;
DFS[16'h11A3] = 8'h00;
DFS[16'h11A4] = 8'h20;
DFS[16'h11A5] = 8'hE1;
DFS[16'h11A6] = 8'h83;
DFS[16'h11A7] = 8'h4C;
DFS[16'h11A8] = 8'hB0;
DFS[16'h11A9] = 8'h91;
DFS[16'h11AA] = 8'h20;
DFS[16'h11AB] = 8'hE1;
DFS[16'h11AC] = 8'h83;
DFS[16'h11AD] = 8'h20;
DFS[16'h11AE] = 8'hA5;
DFS[16'h11AF] = 8'h90;
DFS[16'h11B0] = 8'h48;
DFS[16'h11B1] = 8'hB9;
DFS[16'h11B2] = 8'h0C;
DFS[16'h11B3] = 8'h11;
DFS[16'h11B4] = 8'h30;
DFS[16'h11B5] = 8'hE0;
DFS[16'h11B6] = 8'hB9;
DFS[16'h11B7] = 8'h0E;
DFS[16'h11B8] = 8'h11;
DFS[16'h11B9] = 8'h30;
DFS[16'h11BA] = 8'hD8;
DFS[16'h11BB] = 8'h20;
DFS[16'h11BC] = 8'h83;
DFS[16'h11BD] = 8'h8E;
DFS[16'h11BE] = 8'h98;
DFS[16'h11BF] = 8'h18;
DFS[16'h11C0] = 8'h69;
DFS[16'h11C1] = 8'h04;
DFS[16'h11C2] = 8'h20;
DFS[16'h11C3] = 8'hF8;
DFS[16'h11C4] = 8'h92;
DFS[16'h11C5] = 8'hD0;
DFS[16'h11C6] = 8'h76;
DFS[16'h11C7] = 8'h20;
DFS[16'h11C8] = 8'h58;
DFS[16'h11C9] = 8'h8E;
DFS[16'h11CA] = 8'hAE;
DFS[16'h11CB] = 8'hC4;
DFS[16'h11CC] = 8'h10;
DFS[16'h11CD] = 8'h38;
DFS[16'h11CE] = 8'hBD;
DFS[16'h11CF] = 8'h07;
DFS[16'h11D0] = 8'h0F;
DFS[16'h11D1] = 8'hFD;
DFS[16'h11D2] = 8'h0F;
DFS[16'h11D3] = 8'h0F;
DFS[16'h11D4] = 8'h48;
DFS[16'h11D5] = 8'hBD;
DFS[16'h11D6] = 8'h06;
DFS[16'h11D7] = 8'h0F;
DFS[16'h11D8] = 8'hFD;
DFS[16'h11D9] = 8'h0E;
DFS[16'h11DA] = 8'h0F;
DFS[16'h11DB] = 8'h29;
DFS[16'h11DC] = 8'h03;
DFS[16'h11DD] = 8'h8D;
DFS[16'h11DE] = 8'hC3;
DFS[16'h11DF] = 8'h10;
DFS[16'h11E0] = 8'h0A;
DFS[16'h11E1] = 8'h0A;
DFS[16'h11E2] = 8'h0A;
DFS[16'h11E3] = 8'h0A;
DFS[16'h11E4] = 8'h5D;
DFS[16'h11E5] = 8'h0E;
DFS[16'h11E6] = 8'h0F;
DFS[16'h11E7] = 8'h29;
DFS[16'h11E8] = 8'h30;
DFS[16'h11E9] = 8'h5D;
DFS[16'h11EA] = 8'h0E;
DFS[16'h11EB] = 8'h0F;
DFS[16'h11EC] = 8'h9D;
DFS[16'h11ED] = 8'h0E;
DFS[16'h11EE] = 8'h0F;
DFS[16'h11EF] = 8'hAD;
DFS[16'h11F0] = 8'hC3;
DFS[16'h11F1] = 8'h10;
DFS[16'h11F2] = 8'hD9;
DFS[16'h11F3] = 8'h1A;
DFS[16'h11F4] = 8'h11;
DFS[16'h11F5] = 8'hD0;
DFS[16'h11F6] = 8'h2B;
DFS[16'h11F7] = 8'h68;
DFS[16'h11F8] = 8'hD9;
DFS[16'h11F9] = 8'h19;
DFS[16'h11FA] = 8'h11;
DFS[16'h11FB] = 8'hD0;
DFS[16'h11FC] = 8'h26;
DFS[16'h11FD] = 8'h84;
DFS[16'h11FE] = 8'hB4;
DFS[16'h11FF] = 8'h20;
DFS[16'h1200] = 8'h20;
DFS[16'h1201] = 8'h99;
DFS[16'h1202] = 8'h20;
DFS[16'h1203] = 8'h76;
DFS[16'h1204] = 8'h90;
DFS[16'h1205] = 8'hC4;
DFS[16'h1206] = 8'hB4;
DFS[16'h1207] = 8'hD0;
DFS[16'h1208] = 8'h03;
DFS[16'h1209] = 8'h20;
DFS[16'h120A] = 8'h11;
DFS[16'h120B] = 8'h99;
DFS[16'h120C] = 8'hA4;
DFS[16'h120D] = 8'hB4;
DFS[16'h120E] = 8'h20;
DFS[16'h120F] = 8'h05;
DFS[16'h1210] = 8'h8E;
DFS[16'h1211] = 8'h20;
DFS[16'h1212] = 8'h33;
DFS[16'h1213] = 8'h80;
DFS[16'h1214] = 8'hBF;
DFS[16'h1215] = 8'h43;
DFS[16'h1216] = 8'h61;
DFS[16'h1217] = 8'h6E;
DFS[16'h1218] = 8'h27;
DFS[16'h1219] = 8'h74;
DFS[16'h121A] = 8'h20;
DFS[16'h121B] = 8'h65;
DFS[16'h121C] = 8'h78;
DFS[16'h121D] = 8'h74;
DFS[16'h121E] = 8'h65;
DFS[16'h121F] = 8'h6E;
DFS[16'h1220] = 8'h64;
DFS[16'h1221] = 8'h00;
DFS[16'h1222] = 8'h68;
DFS[16'h1223] = 8'h9D;
DFS[16'h1224] = 8'h0D;
DFS[16'h1225] = 8'h0F;
DFS[16'h1226] = 8'h99;
DFS[16'h1227] = 8'h19;
DFS[16'h1228] = 8'h11;
DFS[16'h1229] = 8'hAD;
DFS[16'h122A] = 8'hC3;
DFS[16'h122B] = 8'h10;
DFS[16'h122C] = 8'h99;
DFS[16'h122D] = 8'h1A;
DFS[16'h122E] = 8'h11;
DFS[16'h122F] = 8'hA9;
DFS[16'h1230] = 8'h00;
DFS[16'h1231] = 8'h9D;
DFS[16'h1232] = 8'h0C;
DFS[16'h1233] = 8'h0F;
DFS[16'h1234] = 8'h20;
DFS[16'h1235] = 8'hB4;
DFS[16'h1236] = 8'h8A;
DFS[16'h1237] = 8'hEA;
DFS[16'h1238] = 8'hEA;
DFS[16'h1239] = 8'hEA;
DFS[16'h123A] = 8'hAC;
DFS[16'h123B] = 8'hC2;
DFS[16'h123C] = 8'h10;
DFS[16'h123D] = 8'hB9;
DFS[16'h123E] = 8'h17;
DFS[16'h123F] = 8'h11;
DFS[16'h1240] = 8'h30;
DFS[16'h1241] = 8'h17;
DFS[16'h1242] = 8'h20;
DFS[16'h1243] = 8'h4B;
DFS[16'h1244] = 8'h91;
DFS[16'h1245] = 8'hB9;
DFS[16'h1246] = 8'h14;
DFS[16'h1247] = 8'h11;
DFS[16'h1248] = 8'hD0;
DFS[16'h1249] = 8'h0B;
DFS[16'h124A] = 8'h98;
DFS[16'h124B] = 8'h20;
DFS[16'h124C] = 8'hF8;
DFS[16'h124D] = 8'h92;
DFS[16'h124E] = 8'hD0;
DFS[16'h124F] = 8'h05;
DFS[16'h1250] = 8'h20;
DFS[16'h1251] = 8'h21;
DFS[16'h1252] = 8'h91;
DFS[16'h1253] = 8'hD0;
DFS[16'h1254] = 8'h04;
DFS[16'h1255] = 8'h38;
DFS[16'h1256] = 8'h20;
DFS[16'h1257] = 8'h53;
DFS[16'h1258] = 8'h91;
DFS[16'h1259] = 8'hB9;
DFS[16'h125A] = 8'h10;
DFS[16'h125B] = 8'h11;
DFS[16'h125C] = 8'h85;
DFS[16'h125D] = 8'hBC;
DFS[16'h125E] = 8'hB9;
DFS[16'h125F] = 8'h13;
DFS[16'h1260] = 8'h11;
DFS[16'h1261] = 8'h85;
DFS[16'h1262] = 8'hBD;
DFS[16'h1263] = 8'h68;
DFS[16'h1264] = 8'hA0;
DFS[16'h1265] = 8'h00;
DFS[16'h1266] = 8'h91;
DFS[16'h1267] = 8'hBC;
DFS[16'h1268] = 8'hAC;
DFS[16'h1269] = 8'hC2;
DFS[16'h126A] = 8'h10;
DFS[16'h126B] = 8'hA9;
DFS[16'h126C] = 8'h40;
DFS[16'h126D] = 8'h20;
DFS[16'h126E] = 8'h3C;
DFS[16'h126F] = 8'h91;
DFS[16'h1270] = 8'hE6;
DFS[16'h1271] = 8'hBC;
DFS[16'h1272] = 8'hA5;
DFS[16'h1273] = 8'hBC;
DFS[16'h1274] = 8'h99;
DFS[16'h1275] = 8'h10;
DFS[16'h1276] = 8'h11;
DFS[16'h1277] = 8'hD0;
DFS[16'h1278] = 8'h13;
DFS[16'h1279] = 8'h20;
DFS[16'h127A] = 8'h41;
DFS[16'h127B] = 8'h91;
DFS[16'h127C] = 8'hB9;
DFS[16'h127D] = 8'h11;
DFS[16'h127E] = 8'h11;
DFS[16'h127F] = 8'h69;
DFS[16'h1280] = 8'h01;
DFS[16'h1281] = 8'h99;
DFS[16'h1282] = 8'h11;
DFS[16'h1283] = 8'h11;
DFS[16'h1284] = 8'hB9;
DFS[16'h1285] = 8'h12;
DFS[16'h1286] = 8'h11;
DFS[16'h1287] = 8'h69;
DFS[16'h1288] = 8'h00;
DFS[16'h1289] = 8'h99;
DFS[16'h128A] = 8'h12;
DFS[16'h128B] = 8'h11;
DFS[16'h128C] = 8'h98;
DFS[16'h128D] = 8'h20;
DFS[16'h128E] = 8'hF8;
DFS[16'h128F] = 8'h92;
DFS[16'h1290] = 8'h90;
DFS[16'h1291] = 8'h14;
DFS[16'h1292] = 8'hA9;
DFS[16'h1293] = 8'h20;
DFS[16'h1294] = 8'h20;
DFS[16'h1295] = 8'h3C;
DFS[16'h1296] = 8'h91;
DFS[16'h1297] = 8'hA2;
DFS[16'h1298] = 8'h02;
DFS[16'h1299] = 8'hB9;
DFS[16'h129A] = 8'h10;
DFS[16'h129B] = 8'h11;
DFS[16'h129C] = 8'h99;
DFS[16'h129D] = 8'h14;
DFS[16'h129E] = 8'h11;
DFS[16'h129F] = 8'hC8;
DFS[16'h12A0] = 8'hCA;
DFS[16'h12A1] = 8'h10;
DFS[16'h12A2] = 8'hF6;
DFS[16'h12A3] = 8'h88;
DFS[16'h12A4] = 8'h88;
DFS[16'h12A5] = 8'h88;
DFS[16'h12A6] = 8'h60;
DFS[16'h12A7] = 8'h20;
DFS[16'h12A8] = 8'hE1;
DFS[16'h12A9] = 8'h83;
DFS[16'h12AA] = 8'h20;
DFS[16'h12AB] = 8'hA5;
DFS[16'h12AC] = 8'h90;
DFS[16'h12AD] = 8'h20;
DFS[16'h12AE] = 8'h5E;
DFS[16'h12AF] = 8'hA1;
DFS[16'h12B0] = 8'hEA;
DFS[16'h12B1] = 8'hEA;
DFS[16'h12B2] = 8'hEA;
DFS[16'h12B3] = 8'hEA;
DFS[16'h12B4] = 8'hEA;
DFS[16'h12B5] = 8'hEA;
DFS[16'h12B6] = 8'h20;
DFS[16'h12B7] = 8'h10;
DFS[16'h12B8] = 8'h93;
DFS[16'h12B9] = 8'hB0;
DFS[16'h12BA] = 8'h08;
DFS[16'h12BB] = 8'hA9;
DFS[16'h12BC] = 8'h00;
DFS[16'h12BD] = 8'h20;
DFS[16'h12BE] = 8'hA4;
DFS[16'h12BF] = 8'h91;
DFS[16'h12C0] = 8'h4C;
DFS[16'h12C1] = 8'hB6;
DFS[16'h12C2] = 8'h92;
DFS[16'h12C3] = 8'hB5;
DFS[16'h12C4] = 8'h00;
DFS[16'h12C5] = 8'h99;
DFS[16'h12C6] = 8'h10;
DFS[16'h12C7] = 8'h11;
DFS[16'h12C8] = 8'hB5;
DFS[16'h12C9] = 8'h01;
DFS[16'h12CA] = 8'h99;
DFS[16'h12CB] = 8'h11;
DFS[16'h12CC] = 8'h11;
DFS[16'h12CD] = 8'hB5;
DFS[16'h12CE] = 8'h02;
DFS[16'h12CF] = 8'h99;
DFS[16'h12D0] = 8'h12;
DFS[16'h12D1] = 8'h11;
DFS[16'h12D2] = 8'hA9;
DFS[16'h12D3] = 8'h6F;
DFS[16'h12D4] = 8'h20;
DFS[16'h12D5] = 8'h43;
DFS[16'h12D6] = 8'h91;
DFS[16'h12D7] = 8'hB9;
DFS[16'h12D8] = 8'h0F;
DFS[16'h12D9] = 8'h11;
DFS[16'h12DA] = 8'h79;
DFS[16'h12DB] = 8'h11;
DFS[16'h12DC] = 8'h11;
DFS[16'h12DD] = 8'h8D;
DFS[16'h12DE] = 8'hC5;
DFS[16'h12DF] = 8'h10;
DFS[16'h12E0] = 8'hB9;
DFS[16'h12E1] = 8'h0D;
DFS[16'h12E2] = 8'h11;
DFS[16'h12E3] = 8'h29;
DFS[16'h12E4] = 8'h03;
DFS[16'h12E5] = 8'h79;
DFS[16'h12E6] = 8'h12;
DFS[16'h12E7] = 8'h11;
DFS[16'h12E8] = 8'hD9;
DFS[16'h12E9] = 8'h1D;
DFS[16'h12EA] = 8'h11;
DFS[16'h12EB] = 8'hD0;
DFS[16'h12EC] = 8'hB9;
DFS[16'h12ED] = 8'hAD;
DFS[16'h12EE] = 8'hC5;
DFS[16'h12EF] = 8'h10;
DFS[16'h12F0] = 8'hD9;
DFS[16'h12F1] = 8'h1C;
DFS[16'h12F2] = 8'h11;
DFS[16'h12F3] = 8'hD0;
DFS[16'h12F4] = 8'hB1;
DFS[16'h12F5] = 8'h4C;
DFS[16'h12F6] = 8'h3A;
DFS[16'h12F7] = 8'h91;
DFS[16'h12F8] = 8'hAA;
DFS[16'h12F9] = 8'hB9;
DFS[16'h12FA] = 8'h12;
DFS[16'h12FB] = 8'h11;
DFS[16'h12FC] = 8'hDD;
DFS[16'h12FD] = 8'h16;
DFS[16'h12FE] = 8'h11;
DFS[16'h12FF] = 8'hD0;
DFS[16'h1300] = 8'h0E;
DFS[16'h1301] = 8'hB9;
DFS[16'h1302] = 8'h11;
DFS[16'h1303] = 8'h11;
DFS[16'h1304] = 8'hDD;
DFS[16'h1305] = 8'h15;
DFS[16'h1306] = 8'h11;
DFS[16'h1307] = 8'hD0;
DFS[16'h1308] = 8'h06;
DFS[16'h1309] = 8'hB9;
DFS[16'h130A] = 8'h10;
DFS[16'h130B] = 8'h11;
DFS[16'h130C] = 8'hDD;
DFS[16'h130D] = 8'h14;
DFS[16'h130E] = 8'h11;
DFS[16'h130F] = 8'h60;
DFS[16'h1310] = 8'hB9;
DFS[16'h1311] = 8'h14;
DFS[16'h1312] = 8'h11;
DFS[16'h1313] = 8'hD5;
DFS[16'h1314] = 8'h00;
DFS[16'h1315] = 8'hB9;
DFS[16'h1316] = 8'h15;
DFS[16'h1317] = 8'h11;
DFS[16'h1318] = 8'hF5;
DFS[16'h1319] = 8'h01;
DFS[16'h131A] = 8'hB9;
DFS[16'h131B] = 8'h16;
DFS[16'h131C] = 8'h11;
DFS[16'h131D] = 8'hF5;
DFS[16'h131E] = 8'h02;
DFS[16'h131F] = 8'h60;
DFS[16'h1320] = 8'hA5;
DFS[16'h1321] = 8'hB3;
DFS[16'h1322] = 8'h48;
DFS[16'h1323] = 8'hA9;
DFS[16'h1324] = 8'hFF;
DFS[16'h1325] = 8'h8D;
DFS[16'h1326] = 8'hDE;
DFS[16'h1327] = 8'h10;
DFS[16'h1328] = 8'h20;
DFS[16'h1329] = 8'h65;
DFS[16'h132A] = 8'h80;
DFS[16'h132B] = 8'h53;
DFS[16'h132C] = 8'h75;
DFS[16'h132D] = 8'h70;
DFS[16'h132E] = 8'h65;
DFS[16'h132F] = 8'h72;
DFS[16'h1330] = 8'h20;
DFS[16'h1331] = 8'h4D;
DFS[16'h1332] = 8'h4D;
DFS[16'h1333] = 8'h43;
DFS[16'h1334] = 8'h0D;
DFS[16'h1335] = 8'h0D;
DFS[16'h1336] = 8'h90;
DFS[16'h1337] = 8'h03;
DFS[16'h1338] = 8'h4C;
DFS[16'h1339] = 8'h55;
DFS[16'h133A] = 8'hA1;
DFS[16'h133B] = 8'hA9;
DFS[16'h133C] = 8'h00;
DFS[16'h133D] = 8'hBA;
DFS[16'h133E] = 8'h9D;
DFS[16'h133F] = 8'h06;
DFS[16'h1340] = 8'h01;
DFS[16'h1341] = 8'hA9;
DFS[16'h1342] = 8'h06;
DFS[16'h1343] = 8'h20;
DFS[16'h1344] = 8'h15;
DFS[16'h1345] = 8'h80;
DFS[16'h1346] = 8'hA2;
DFS[16'h1347] = 8'h0D;
DFS[16'h1348] = 8'hBD;
DFS[16'h1349] = 8'h49;
DFS[16'h134A] = 8'h99;
DFS[16'h134B] = 8'h9D;
DFS[16'h134C] = 8'h12;
DFS[16'h134D] = 8'h02;
DFS[16'h134E] = 8'hCA;
DFS[16'h134F] = 8'h10;
DFS[16'h1350] = 8'hF7;
DFS[16'h1351] = 8'h20;
DFS[16'h1352] = 8'h28;
DFS[16'h1353] = 8'h99;
DFS[16'h1354] = 8'h84;
DFS[16'h1355] = 8'hB1;
DFS[16'h1356] = 8'h86;
DFS[16'h1357] = 8'hB0;
DFS[16'h1358] = 8'hA2;
DFS[16'h1359] = 8'h07;
DFS[16'h135A] = 8'hA0;
DFS[16'h135B] = 8'h1B;
DFS[16'h135C] = 8'hB9;
DFS[16'h135D] = 8'h3C;
DFS[16'h135E] = 8'h99;
DFS[16'h135F] = 8'h91;
DFS[16'h1360] = 8'hB0;
DFS[16'h1361] = 8'hC8;
DFS[16'h1362] = 8'hB9;
DFS[16'h1363] = 8'h3C;
DFS[16'h1364] = 8'h99;
DFS[16'h1365] = 8'h91;
DFS[16'h1366] = 8'hB0;
DFS[16'h1367] = 8'hC8;
DFS[16'h1368] = 8'hA5;
DFS[16'h1369] = 8'hF4;
DFS[16'h136A] = 8'h91;
DFS[16'h136B] = 8'hB0;
DFS[16'h136C] = 8'hC8;
DFS[16'h136D] = 8'hCA;
DFS[16'h136E] = 8'hD0;
DFS[16'h136F] = 8'hEC;
DFS[16'h1370] = 8'h86;
DFS[16'h1371] = 8'hCF;
DFS[16'h1372] = 8'h8C;
DFS[16'h1373] = 8'h82;
DFS[16'h1374] = 8'h10;
DFS[16'h1375] = 8'hA2;
DFS[16'h1376] = 8'h0F;
DFS[16'h1377] = 8'h20;
DFS[16'h1378] = 8'h2C;
DFS[16'h1379] = 8'h99;
DFS[16'h137A] = 8'h20;
DFS[16'h137B] = 8'h9E;
DFS[16'h137C] = 8'h98;
DFS[16'h137D] = 8'hA0;
DFS[16'h137E] = 8'hD4;
DFS[16'h137F] = 8'hB1;
DFS[16'h1380] = 8'hB0;
DFS[16'h1381] = 8'h10;
DFS[16'h1382] = 8'h2F;
DFS[16'h1383] = 8'hA0;
DFS[16'h1384] = 8'hD5;
DFS[16'h1385] = 8'hB1;
DFS[16'h1386] = 8'hB0;
DFS[16'h1387] = 8'h30;
DFS[16'h1388] = 8'h27;
DFS[16'h1389] = 8'h20;
DFS[16'h138A] = 8'h8F;
DFS[16'h138B] = 8'h98;
DFS[16'h138C] = 8'hA0;
DFS[16'h138D] = 8'h00;
DFS[16'h138E] = 8'hB1;
DFS[16'h138F] = 8'hB0;
DFS[16'h1390] = 8'hC0;
DFS[16'h1391] = 8'hC0;
DFS[16'h1392] = 8'h90;
DFS[16'h1393] = 8'h05;
DFS[16'h1394] = 8'h99;
DFS[16'h1395] = 8'h00;
DFS[16'h1396] = 8'h10;
DFS[16'h1397] = 8'hB0;
DFS[16'h1398] = 8'h03;
DFS[16'h1399] = 8'h99;
DFS[16'h139A] = 8'h00;
DFS[16'h139B] = 8'h11;
DFS[16'h139C] = 8'h88;
DFS[16'h139D] = 8'hD0;
DFS[16'h139E] = 8'hEF;
DFS[16'h139F] = 8'hA9;
DFS[16'h13A0] = 8'hA0;
DFS[16'h13A1] = 8'hA8;
DFS[16'h13A2] = 8'h48;
DFS[16'h13A3] = 8'hA9;
DFS[16'h13A4] = 8'h3F;
DFS[16'h13A5] = 8'h20;
DFS[16'h13A6] = 8'h43;
DFS[16'h13A7] = 8'h91;
DFS[16'h13A8] = 8'h68;
DFS[16'h13A9] = 8'h99;
DFS[16'h13AA] = 8'h1D;
DFS[16'h13AB] = 8'h11;
DFS[16'h13AC] = 8'hE9;
DFS[16'h13AD] = 8'h1F;
DFS[16'h13AE] = 8'hD0;
DFS[16'h13AF] = 8'hF1;
DFS[16'h13B0] = 8'h68;
DFS[16'h13B1] = 8'h60;
DFS[16'h13B2] = 8'hA9;
DFS[16'h13B3] = 8'hFF;
DFS[16'h13B4] = 8'h91;
DFS[16'h13B5] = 8'hB0;
DFS[16'h13B6] = 8'h8D;
DFS[16'h13B7] = 8'hD4;
DFS[16'h13B8] = 8'h10;
DFS[16'h13B9] = 8'h20;
DFS[16'h13BA] = 8'h8F;
DFS[16'h13BB] = 8'h98;
DFS[16'h13BC] = 8'h20;
DFS[16'h13BD] = 8'h24;
DFS[16'h13BE] = 8'h99;
DFS[16'h13BF] = 8'h8A;
DFS[16'h13C0] = 8'h49;
DFS[16'h13C1] = 8'hFF;
DFS[16'h13C2] = 8'h8D;
DFS[16'h13C3] = 8'hD7;
DFS[16'h13C4] = 8'h10;
DFS[16'h13C5] = 8'hA9;
DFS[16'h13C6] = 8'h24;
DFS[16'h13C7] = 8'h8D;
DFS[16'h13C8] = 8'hCA;
DFS[16'h13C9] = 8'h10;
DFS[16'h13CA] = 8'h8D;
DFS[16'h13CB] = 8'hCC;
DFS[16'h13CC] = 8'h10;
DFS[16'h13CD] = 8'hA0;
DFS[16'h13CE] = 8'h00;
DFS[16'h13CF] = 8'h8C;
DFS[16'h13D0] = 8'hCB;
DFS[16'h13D1] = 8'h10;
DFS[16'h13D2] = 8'h8C;
DFS[16'h13D3] = 8'hCD;
DFS[16'h13D4] = 8'h10;
DFS[16'h13D5] = 8'hA0;
DFS[16'h13D6] = 8'h00;
DFS[16'h13D7] = 8'h8C;
DFS[16'h13D8] = 8'hC0;
DFS[16'h13D9] = 8'h10;
DFS[16'h13DA] = 8'h8C;
DFS[16'h13DB] = 8'hC9;
DFS[16'h13DC] = 8'h10;
DFS[16'h13DD] = 8'h88;
DFS[16'h13DE] = 8'h8C;
DFS[16'h13DF] = 8'hC8;
DFS[16'h13E0] = 8'h10;
DFS[16'h13E1] = 8'h8C;
DFS[16'h13E2] = 8'hC7;
DFS[16'h13E3] = 8'h10;
DFS[16'h13E4] = 8'h8C;
DFS[16'h13E5] = 8'hDE;
DFS[16'h13E6] = 8'h10;
DFS[16'h13E7] = 8'h20;
DFS[16'h13E8] = 8'h0A;
DFS[16'h13E9] = 8'hAD;
DFS[16'h13EA] = 8'h4C;
DFS[16'h13EB] = 8'h04;
DFS[16'h13EC] = 8'h94;
DFS[16'h13ED] = 8'h00;
DFS[16'h13EE] = 8'h00;
DFS[16'h13EF] = 8'h00;
DFS[16'h13F0] = 8'h00;
DFS[16'h13F1] = 8'h00;
DFS[16'h13F2] = 8'h00;
DFS[16'h13F3] = 8'h00;
DFS[16'h13F4] = 8'h00;
DFS[16'h13F5] = 8'h00;
DFS[16'h13F6] = 8'h00;
DFS[16'h13F7] = 8'h00;
DFS[16'h13F8] = 8'h00;
DFS[16'h13F9] = 8'h00;
DFS[16'h13FA] = 8'h00;
DFS[16'h13FB] = 8'h00;
DFS[16'h13FC] = 8'h00;
DFS[16'h13FD] = 8'h00;
DFS[16'h13FE] = 8'h00;
DFS[16'h13FF] = 8'h00;
DFS[16'h1400] = 8'h00;
DFS[16'h1401] = 8'h00;
DFS[16'h1402] = 8'h00;
DFS[16'h1403] = 8'h00;
DFS[16'h1404] = 8'h68;
DFS[16'h1405] = 8'hD0;
DFS[16'h1406] = 8'h34;
DFS[16'h1407] = 8'h20;
DFS[16'h1408] = 8'h4D;
DFS[16'h1409] = 8'hAB;
DFS[16'h140A] = 8'hA0;
DFS[16'h140B] = 8'h00;
DFS[16'h140C] = 8'hA2;
DFS[16'h140D] = 8'h00;
DFS[16'h140E] = 8'hAD;
DFS[16'h140F] = 8'h06;
DFS[16'h1410] = 8'h0F;
DFS[16'h1411] = 8'h20;
DFS[16'h1412] = 8'h05;
DFS[16'h1413] = 8'h82;
DFS[16'h1414] = 8'hF0;
DFS[16'h1415] = 8'h25;
DFS[16'h1416] = 8'h48;
DFS[16'h1417] = 8'hA2;
DFS[16'h1418] = 8'h43;
DFS[16'h1419] = 8'hA0;
DFS[16'h141A] = 8'h99;
DFS[16'h141B] = 8'h20;
DFS[16'h141C] = 8'hB8;
DFS[16'h141D] = 8'h86;
DFS[16'h141E] = 8'h20;
DFS[16'h141F] = 8'hFE;
DFS[16'h1420] = 8'h80;
DFS[16'h1421] = 8'h20;
DFS[16'h1422] = 8'h96;
DFS[16'h1423] = 8'h82;
DFS[16'h1424] = 8'h68;
DFS[16'h1425] = 8'hB0;
DFS[16'h1426] = 8'h15;
DFS[16'h1427] = 8'h20;
DFS[16'h1428] = 8'h65;
DFS[16'h1429] = 8'h80;
DFS[16'h142A] = 8'h46;
DFS[16'h142B] = 8'h69;
DFS[16'h142C] = 8'h6C;
DFS[16'h142D] = 8'h65;
DFS[16'h142E] = 8'h20;
DFS[16'h142F] = 8'h6E;
DFS[16'h1430] = 8'h6F;
DFS[16'h1431] = 8'h74;
DFS[16'h1432] = 8'h20;
DFS[16'h1433] = 8'h66;
DFS[16'h1434] = 8'h6F;
DFS[16'h1435] = 8'h75;
DFS[16'h1436] = 8'h6E;
DFS[16'h1437] = 8'h64;
DFS[16'h1438] = 8'h0D;
DFS[16'h1439] = 8'h0D;
DFS[16'h143A] = 8'hEA;
DFS[16'h143B] = 8'h60;
DFS[16'h143C] = 8'hC9;
DFS[16'h143D] = 8'h02;
DFS[16'h143E] = 8'h90;
DFS[16'h143F] = 8'h0E;
DFS[16'h1440] = 8'hF0;
DFS[16'h1441] = 8'h06;
DFS[16'h1442] = 8'hA2;
DFS[16'h1443] = 8'h41;
DFS[16'h1444] = 8'hA0;
DFS[16'h1445] = 8'h99;
DFS[16'h1446] = 8'hD0;
DFS[16'h1447] = 8'h0A;
DFS[16'h1448] = 8'hA2;
DFS[16'h1449] = 8'h43;
DFS[16'h144A] = 8'hA0;
DFS[16'h144B] = 8'h99;
DFS[16'h144C] = 8'hD0;
DFS[16'h144D] = 8'h04;
DFS[16'h144E] = 8'hA2;
DFS[16'h144F] = 8'h39;
DFS[16'h1450] = 8'hA0;
DFS[16'h1451] = 8'h99;
DFS[16'h1452] = 8'h4C;
DFS[16'h1453] = 8'hF7;
DFS[16'h1454] = 8'hFF;
DFS[16'h1455] = 8'hC9;
DFS[16'h1456] = 8'h01;
DFS[16'h1457] = 8'hD0;
DFS[16'h1458] = 8'h07;
DFS[16'h1459] = 8'hC0;
DFS[16'h145A] = 8'h17;
DFS[16'h145B] = 8'hB0;
DFS[16'h145C] = 8'h02;
DFS[16'h145D] = 8'hA0;
DFS[16'h145E] = 8'h17;
DFS[16'h145F] = 8'h60;
DFS[16'h1460] = 8'hC9;
DFS[16'h1461] = 8'h02;
DFS[16'h1462] = 8'hD0;
DFS[16'h1463] = 8'h1A;
DFS[16'h1464] = 8'h48;
DFS[16'h1465] = 8'h98;
DFS[16'h1466] = 8'h18;
DFS[16'h1467] = 8'h85;
DFS[16'h1468] = 8'hB1;
DFS[16'h1469] = 8'h9D;
DFS[16'h146A] = 8'hF0;
DFS[16'h146B] = 8'h0D;
DFS[16'h146C] = 8'h69;
DFS[16'h146D] = 8'h02;
DFS[16'h146E] = 8'h48;
DFS[16'h146F] = 8'hA9;
DFS[16'h1470] = 8'h00;
DFS[16'h1471] = 8'h85;
DFS[16'h1472] = 8'hB0;
DFS[16'h1473] = 8'hA0;
DFS[16'h1474] = 8'hD4;
DFS[16'h1475] = 8'h91;
DFS[16'h1476] = 8'hB0;
DFS[16'h1477] = 8'hC8;
DFS[16'h1478] = 8'h91;
DFS[16'h1479] = 8'hB0;
DFS[16'h147A] = 8'h68;
DFS[16'h147B] = 8'hA8;
DFS[16'h147C] = 8'h68;
DFS[16'h147D] = 8'h60;
DFS[16'h147E] = 8'hC9;
DFS[16'h147F] = 8'h03;
DFS[16'h1480] = 8'hD0;
DFS[16'h1481] = 8'h19;
DFS[16'h1482] = 8'h84;
DFS[16'h1483] = 8'hB3;
DFS[16'h1484] = 8'h20;
DFS[16'h1485] = 8'hE1;
DFS[16'h1486] = 8'h83;
DFS[16'h1487] = 8'h4C;
DFS[16'h1488] = 8'hF7;
DFS[16'h1489] = 8'hA7;
DFS[16'h148A] = 8'hF4;
DFS[16'h148B] = 8'hFF;
DFS[16'h148C] = 8'h8A;
DFS[16'h148D] = 8'h30;
DFS[16'h148E] = 8'h09;
DFS[16'h148F] = 8'hC9;
DFS[16'h1490] = 8'h32;
DFS[16'h1491] = 8'hD0;
DFS[16'h1492] = 8'hEA;
DFS[16'h1493] = 8'hA9;
DFS[16'h1494] = 8'h78;
DFS[16'h1495] = 8'h20;
DFS[16'h1496] = 8'hF4;
DFS[16'h1497] = 8'hFF;
DFS[16'h1498] = 8'h4C;
DFS[16'h1499] = 8'h20;
DFS[16'h149A] = 8'h93;
DFS[16'h149B] = 8'hC9;
DFS[16'h149C] = 8'h04;
DFS[16'h149D] = 8'hD0;
DFS[16'h149E] = 8'h08;
DFS[16'h149F] = 8'h20;
DFS[16'h14A0] = 8'hE1;
DFS[16'h14A1] = 8'h83;
DFS[16'h14A2] = 8'hA2;
DFS[16'h14A3] = 8'h72;
DFS[16'h14A4] = 8'h4C;
DFS[16'h14A5] = 8'h71;
DFS[16'h14A6] = 8'h86;
DFS[16'h14A7] = 8'hC9;
DFS[16'h14A8] = 8'h09;
DFS[16'h14A9] = 8'hD0;
DFS[16'h14AA] = 8'h12;
DFS[16'h14AB] = 8'h20;
DFS[16'h14AC] = 8'hE1;
DFS[16'h14AD] = 8'h83;
DFS[16'h14AE] = 8'h4C;
DFS[16'h14AF] = 8'h94;
DFS[16'h14B0] = 8'hAF;
DFS[16'h14B1] = 8'hA0;
DFS[16'h14B2] = 8'hC9;
DFS[16'h14B3] = 8'h0D;
DFS[16'h14B4] = 8'hD0;
DFS[16'h14B5] = 8'hEE;
DFS[16'h14B6] = 8'h98;
DFS[16'h14B7] = 8'hE8;
DFS[16'h14B8] = 8'hA0;
DFS[16'h14B9] = 8'h02;
DFS[16'h14BA] = 8'h4C;
DFS[16'h14BB] = 8'hCB;
DFS[16'h14BC] = 8'h99;
DFS[16'h14BD] = 8'hC9;
DFS[16'h14BE] = 8'h0A;
DFS[16'h14BF] = 8'hD0;
DFS[16'h14C0] = 8'h29;
DFS[16'h14C1] = 8'h20;
DFS[16'h14C2] = 8'hE1;
DFS[16'h14C3] = 8'h83;
DFS[16'h14C4] = 8'h20;
DFS[16'h14C5] = 8'h9E;
DFS[16'h14C6] = 8'h98;
DFS[16'h14C7] = 8'hA0;
DFS[16'h14C8] = 8'hD5;
DFS[16'h14C9] = 8'hB1;
DFS[16'h14CA] = 8'hB0;
DFS[16'h14CB] = 8'h10;
DFS[16'h14CC] = 8'h1C;
DFS[16'h14CD] = 8'hA0;
DFS[16'h14CE] = 8'h00;
DFS[16'h14CF] = 8'hC0;
DFS[16'h14D0] = 8'hC0;
DFS[16'h14D1] = 8'h90;
DFS[16'h14D2] = 8'h05;
DFS[16'h14D3] = 8'hB9;
DFS[16'h14D4] = 8'h00;
DFS[16'h14D5] = 8'h10;
DFS[16'h14D6] = 8'hB0;
DFS[16'h14D7] = 8'h03;
DFS[16'h14D8] = 8'hB9;
DFS[16'h14D9] = 8'h00;
DFS[16'h14DA] = 8'h11;
DFS[16'h14DB] = 8'h91;
DFS[16'h14DC] = 8'hB0;
DFS[16'h14DD] = 8'h88;
DFS[16'h14DE] = 8'hD0;
DFS[16'h14DF] = 8'hEF;
DFS[16'h14E0] = 8'h20;
DFS[16'h14E1] = 8'hF2;
DFS[16'h14E2] = 8'h8F;
DFS[16'h14E3] = 8'hA0;
DFS[16'h14E4] = 8'hD5;
DFS[16'h14E5] = 8'hA9;
DFS[16'h14E6] = 8'h00;
DFS[16'h14E7] = 8'h91;
DFS[16'h14E8] = 8'hB0;
DFS[16'h14E9] = 8'h60;
DFS[16'h14EA] = 8'hC9;
DFS[16'h14EB] = 8'h08;
DFS[16'h14EC] = 8'hD0;
DFS[16'h14ED] = 8'h15;
DFS[16'h14EE] = 8'h20;
DFS[16'h14EF] = 8'h11;
DFS[16'h14F0] = 8'h84;
DFS[16'h14F1] = 8'hA4;
DFS[16'h14F2] = 8'hF0;
DFS[16'h14F3] = 8'h84;
DFS[16'h14F4] = 8'hB0;
DFS[16'h14F5] = 8'hA4;
DFS[16'h14F6] = 8'hF1;
DFS[16'h14F7] = 8'h84;
DFS[16'h14F8] = 8'hB1;
DFS[16'h14F9] = 8'hA4;
DFS[16'h14FA] = 8'hEF;
DFS[16'h14FB] = 8'hC0;
DFS[16'h14FC] = 8'h7F;
DFS[16'h14FD] = 8'hD0;
DFS[16'h14FE] = 8'h4C;
DFS[16'h14FF] = 8'h4C;
DFS[16'h1500] = 8'h13;
DFS[16'h1501] = 8'hB9;
DFS[16'h1502] = 8'h00;
DFS[16'h1503] = 8'h4C;
DFS[16'h1504] = 8'hF6;
DFS[16'h1505] = 8'hA0;
DFS[16'h1506] = 8'h00;
DFS[16'h1507] = 8'h00;
DFS[16'h1508] = 8'h00;
DFS[16'h1509] = 8'h00;
DFS[16'h150A] = 8'h00;
DFS[16'h150B] = 8'h00;
DFS[16'h150C] = 8'h00;
DFS[16'h150D] = 8'h00;
DFS[16'h150E] = 8'h00;
DFS[16'h150F] = 8'h00;
DFS[16'h1510] = 8'h00;
DFS[16'h1511] = 8'h00;
DFS[16'h1512] = 8'h00;
DFS[16'h1513] = 8'h00;
DFS[16'h1514] = 8'h00;
DFS[16'h1515] = 8'h00;
DFS[16'h1516] = 8'h00;
DFS[16'h1517] = 8'h00;
DFS[16'h1518] = 8'h00;
DFS[16'h1519] = 8'h00;
DFS[16'h151A] = 8'h00;
DFS[16'h151B] = 8'h00;
DFS[16'h151C] = 8'h00;
DFS[16'h151D] = 8'h00;
DFS[16'h151E] = 8'h00;
DFS[16'h151F] = 8'h00;
DFS[16'h1520] = 8'h00;
DFS[16'h1521] = 8'h00;
DFS[16'h1522] = 8'h00;
DFS[16'h1523] = 8'h00;
DFS[16'h1524] = 8'h00;
DFS[16'h1525] = 8'h00;
DFS[16'h1526] = 8'h00;
DFS[16'h1527] = 8'h00;
DFS[16'h1528] = 8'h00;
DFS[16'h1529] = 8'h00;
DFS[16'h152A] = 8'h00;
DFS[16'h152B] = 8'h00;
DFS[16'h152C] = 8'h00;
DFS[16'h152D] = 8'h00;
DFS[16'h152E] = 8'h00;
DFS[16'h152F] = 8'h00;
DFS[16'h1530] = 8'h00;
DFS[16'h1531] = 8'h00;
DFS[16'h1532] = 8'h00;
DFS[16'h1533] = 8'h00;
DFS[16'h1534] = 8'h00;
DFS[16'h1535] = 8'h00;
DFS[16'h1536] = 8'h00;
DFS[16'h1537] = 8'h00;
DFS[16'h1538] = 8'h00;
DFS[16'h1539] = 8'h00;
DFS[16'h153A] = 8'h00;
DFS[16'h153B] = 8'h00;
DFS[16'h153C] = 8'h00;
DFS[16'h153D] = 8'h00;
DFS[16'h153E] = 8'h00;
DFS[16'h153F] = 8'h00;
DFS[16'h1540] = 8'h00;
DFS[16'h1541] = 8'h00;
DFS[16'h1542] = 8'h00;
DFS[16'h1543] = 8'h00;
DFS[16'h1544] = 8'h00;
DFS[16'h1545] = 8'h00;
DFS[16'h1546] = 8'h00;
DFS[16'h1547] = 8'h00;
DFS[16'h1548] = 8'h00;
DFS[16'h1549] = 8'h00;
DFS[16'h154A] = 8'h00;
DFS[16'h154B] = 8'hC0;
DFS[16'h154C] = 8'h7D;
DFS[16'h154D] = 8'h90;
DFS[16'h154E] = 8'h2B;
DFS[16'h154F] = 8'h20;
DFS[16'h1550] = 8'h4D;
DFS[16'h1551] = 8'h83;
DFS[16'h1552] = 8'h20;
DFS[16'h1553] = 8'h47;
DFS[16'h1554] = 8'h83;
DFS[16'h1555] = 8'hC0;
DFS[16'h1556] = 8'h7E;
DFS[16'h1557] = 8'hF0;
DFS[16'h1558] = 8'h09;
DFS[16'h1559] = 8'hA0;
DFS[16'h155A] = 8'h00;
DFS[16'h155B] = 8'hAD;
DFS[16'h155C] = 8'h04;
DFS[16'h155D] = 8'h0F;
DFS[16'h155E] = 8'h91;
DFS[16'h155F] = 8'hB0;
DFS[16'h1560] = 8'h98;
DFS[16'h1561] = 8'h60;
DFS[16'h1562] = 8'hA9;
DFS[16'h1563] = 8'h00;
DFS[16'h1564] = 8'hA8;
DFS[16'h1565] = 8'h91;
DFS[16'h1566] = 8'hB0;
DFS[16'h1567] = 8'hC8;
DFS[16'h1568] = 8'hAD;
DFS[16'h1569] = 8'h07;
DFS[16'h156A] = 8'h0F;
DFS[16'h156B] = 8'h91;
DFS[16'h156C] = 8'hB0;
DFS[16'h156D] = 8'hC8;
DFS[16'h156E] = 8'hAD;
DFS[16'h156F] = 8'h06;
DFS[16'h1570] = 8'h0F;
DFS[16'h1571] = 8'h29;
DFS[16'h1572] = 8'h03;
DFS[16'h1573] = 8'h91;
DFS[16'h1574] = 8'hB0;
DFS[16'h1575] = 8'hC8;
DFS[16'h1576] = 8'hA9;
DFS[16'h1577] = 8'h00;
DFS[16'h1578] = 8'h91;
DFS[16'h1579] = 8'hB0;
DFS[16'h157A] = 8'h60;
DFS[16'h157B] = 8'h20;
DFS[16'h157C] = 8'h11;
DFS[16'h157D] = 8'h84;
DFS[16'h157E] = 8'h48;
DFS[16'h157F] = 8'h20;
DFS[16'h1580] = 8'h62;
DFS[16'h1581] = 8'h82;
DFS[16'h1582] = 8'h86;
DFS[16'h1583] = 8'hB0;
DFS[16'h1584] = 8'h8E;
DFS[16'h1585] = 8'hDC;
DFS[16'h1586] = 8'h10;
DFS[16'h1587] = 8'h84;
DFS[16'h1588] = 8'hB1;
DFS[16'h1589] = 8'h8C;
DFS[16'h158A] = 8'hDD;
DFS[16'h158B] = 8'h10;
DFS[16'h158C] = 8'hA2;
DFS[16'h158D] = 8'h00;
DFS[16'h158E] = 8'hA0;
DFS[16'h158F] = 8'h00;
DFS[16'h1590] = 8'h20;
DFS[16'h1591] = 8'hEA;
DFS[16'h1592] = 8'h80;
DFS[16'h1593] = 8'h20;
DFS[16'h1594] = 8'hDA;
DFS[16'h1595] = 8'h80;
DFS[16'h1596] = 8'hC0;
DFS[16'h1597] = 8'h12;
DFS[16'h1598] = 8'hD0;
DFS[16'h1599] = 8'hF9;
DFS[16'h159A] = 8'h68;
DFS[16'h159B] = 8'hAA;
DFS[16'h159C] = 8'hE8;
DFS[16'h159D] = 8'hE0;
DFS[16'h159E] = 8'h08;
DFS[16'h159F] = 8'hB0;
DFS[16'h15A0] = 8'h08;
DFS[16'h15A1] = 8'hBD;
DFS[16'h15A2] = 8'h8C;
DFS[16'h15A3] = 8'h99;
DFS[16'h15A4] = 8'h48;
DFS[16'h15A5] = 8'hBD;
DFS[16'h15A6] = 8'h84;
DFS[16'h15A7] = 8'h99;
DFS[16'h15A8] = 8'h48;
DFS[16'h15A9] = 8'h60;
DFS[16'h15AA] = 8'hC9;
DFS[16'h15AB] = 8'h09;
DFS[16'h15AC] = 8'hB0;
DFS[16'h15AD] = 8'hFB;
DFS[16'h15AE] = 8'h86;
DFS[16'h15AF] = 8'hB5;
DFS[16'h15B0] = 8'hAA;
DFS[16'h15B1] = 8'hBD;
DFS[16'h15B2] = 8'h75;
DFS[16'h15B3] = 8'h99;
DFS[16'h15B4] = 8'h48;
DFS[16'h15B5] = 8'hBD;
DFS[16'h15B6] = 8'h6C;
DFS[16'h15B7] = 8'h99;
DFS[16'h15B8] = 8'h48;
DFS[16'h15B9] = 8'h8A;
DFS[16'h15BA] = 8'hA6;
DFS[16'h15BB] = 8'hB5;
DFS[16'h15BC] = 8'h60;
DFS[16'h15BD] = 8'hA9;
DFS[16'h15BE] = 8'hFF;
DFS[16'h15BF] = 8'h95;
DFS[16'h15C0] = 8'h02;
DFS[16'h15C1] = 8'h95;
DFS[16'h15C2] = 8'h03;
DFS[16'h15C3] = 8'hAD;
DFS[16'h15C4] = 8'hDA;
DFS[16'h15C5] = 8'h10;
DFS[16'h15C6] = 8'h95;
DFS[16'h15C7] = 8'h00;
DFS[16'h15C8] = 8'hAD;
DFS[16'h15C9] = 8'hDB;
DFS[16'h15CA] = 8'h10;
DFS[16'h15CB] = 8'h95;
DFS[16'h15CC] = 8'h01;
DFS[16'h15CD] = 8'hA9;
DFS[16'h15CE] = 8'h00;
DFS[16'h15CF] = 8'h60;
DFS[16'h15D0] = 8'hC9;
DFS[16'h15D1] = 8'h09;
DFS[16'h15D2] = 8'hB0;
DFS[16'h15D3] = 8'hFB;
DFS[16'h15D4] = 8'h20;
DFS[16'h15D5] = 8'hE1;
DFS[16'h15D6] = 8'h83;
DFS[16'h15D7] = 8'h8E;
DFS[16'h15D8] = 8'h7D;
DFS[16'h15D9] = 8'h10;
DFS[16'h15DA] = 8'h8C;
DFS[16'h15DB] = 8'h7E;
DFS[16'h15DC] = 8'h10;
DFS[16'h15DD] = 8'hA8;
DFS[16'h15DE] = 8'hBA;
DFS[16'h15DF] = 8'hA9;
DFS[16'h15E0] = 8'h00;
DFS[16'h15E1] = 8'h4C;
DFS[16'h15E2] = 8'hD8;
DFS[16'h15E3] = 8'hA0;
DFS[16'h15E4] = 8'hB9;
DFS[16'h15E5] = 8'hAB;
DFS[16'h15E6] = 8'h99;
DFS[16'h15E7] = 8'h8D;
DFS[16'h15E8] = 8'hD8;
DFS[16'h15E9] = 8'h10;
DFS[16'h15EA] = 8'hB9;
DFS[16'h15EB] = 8'hB4;
DFS[16'h15EC] = 8'h99;
DFS[16'h15ED] = 8'h8D;
DFS[16'h15EE] = 8'hD9;
DFS[16'h15EF] = 8'h10;
DFS[16'h15F0] = 8'hB9;
DFS[16'h15F1] = 8'hBD;
DFS[16'h15F2] = 8'h99;
DFS[16'h15F3] = 8'h4A;
DFS[16'h15F4] = 8'h08;
DFS[16'h15F5] = 8'h4A;
DFS[16'h15F6] = 8'h08;
DFS[16'h15F7] = 8'h8D;
DFS[16'h15F8] = 8'h7F;
DFS[16'h15F9] = 8'h10;
DFS[16'h15FA] = 8'h20;
DFS[16'h15FB] = 8'h56;
DFS[16'h15FC] = 8'h97;
DFS[16'h15FD] = 8'hA0;
DFS[16'h15FE] = 8'h0C;
DFS[16'h15FF] = 8'hB1;
DFS[16'h1600] = 8'hB4;
DFS[16'h1601] = 8'h99;
DFS[16'h1602] = 8'h60;
DFS[16'h1603] = 8'h10;
DFS[16'h1604] = 8'h88;
DFS[16'h1605] = 8'h10;
DFS[16'h1606] = 8'hF8;
DFS[16'h1607] = 8'hAD;
DFS[16'h1608] = 8'h63;
DFS[16'h1609] = 8'h10;
DFS[16'h160A] = 8'h2D;
DFS[16'h160B] = 8'h64;
DFS[16'h160C] = 8'h10;
DFS[16'h160D] = 8'h0D;
DFS[16'h160E] = 8'hD7;
DFS[16'h160F] = 8'h10;
DFS[16'h1610] = 8'h18;
DFS[16'h1611] = 8'h69;
DFS[16'h1612] = 8'h01;
DFS[16'h1613] = 8'h4C;
DFS[16'h1614] = 8'hEB;
DFS[16'h1615] = 8'hA0;
DFS[16'h1616] = 8'hEA;
DFS[16'h1617] = 8'h8D;
DFS[16'h1618] = 8'h81;
DFS[16'h1619] = 8'h10;
DFS[16'h161A] = 8'hAD;
DFS[16'h161B] = 8'h7F;
DFS[16'h161C] = 8'h10;
DFS[16'h161D] = 8'hB0;
DFS[16'h161E] = 8'h07;
DFS[16'h161F] = 8'hA2;
DFS[16'h1620] = 8'h61;
DFS[16'h1621] = 8'hA0;
DFS[16'h1622] = 8'h10;
DFS[16'h1623] = 8'h20;
DFS[16'h1624] = 8'h06;
DFS[16'h1625] = 8'h04;
DFS[16'h1626] = 8'h28;
DFS[16'h1627] = 8'hB0;
DFS[16'h1628] = 8'h04;
DFS[16'h1629] = 8'h28;
DFS[16'h162A] = 8'h6C;
DFS[16'h162B] = 8'hD8;
DFS[16'h162C] = 8'h10;
DFS[16'h162D] = 8'hA2;
DFS[16'h162E] = 8'h03;
DFS[16'h162F] = 8'hBD;
DFS[16'h1630] = 8'h69;
DFS[16'h1631] = 8'h10;
DFS[16'h1632] = 8'h95;
DFS[16'h1633] = 8'hB6;
DFS[16'h1634] = 8'hCA;
DFS[16'h1635] = 8'h10;
DFS[16'h1636] = 8'hF8;
DFS[16'h1637] = 8'hA2;
DFS[16'h1638] = 8'hB6;
DFS[16'h1639] = 8'hAC;
DFS[16'h163A] = 8'h60;
DFS[16'h163B] = 8'h10;
DFS[16'h163C] = 8'hA9;
DFS[16'h163D] = 8'h00;
DFS[16'h163E] = 8'h28;
DFS[16'h163F] = 8'hB0;
DFS[16'h1640] = 8'h03;
DFS[16'h1641] = 8'h20;
DFS[16'h1642] = 8'hA7;
DFS[16'h1643] = 8'h92;
DFS[16'h1644] = 8'h20;
DFS[16'h1645] = 8'h2E;
DFS[16'h1646] = 8'h90;
DFS[16'h1647] = 8'hA2;
DFS[16'h1648] = 8'h03;
DFS[16'h1649] = 8'hB5;
DFS[16'h164A] = 8'hB6;
DFS[16'h164B] = 8'h9D;
DFS[16'h164C] = 8'h69;
DFS[16'h164D] = 8'h10;
DFS[16'h164E] = 8'hCA;
DFS[16'h164F] = 8'h10;
DFS[16'h1650] = 8'hF8;
DFS[16'h1651] = 8'h20;
DFS[16'h1652] = 8'h48;
DFS[16'h1653] = 8'h97;
DFS[16'h1654] = 8'h30;
DFS[16'h1655] = 8'h0D;
DFS[16'h1656] = 8'hAC;
DFS[16'h1657] = 8'h60;
DFS[16'h1658] = 8'h10;
DFS[16'h1659] = 8'h20;
DFS[16'h165A] = 8'h2A;
DFS[16'h165B] = 8'h96;
DFS[16'h165C] = 8'hB0;
DFS[16'h165D] = 8'h0D;
DFS[16'h165E] = 8'hA2;
DFS[16'h165F] = 8'h09;
DFS[16'h1660] = 8'h20;
DFS[16'h1661] = 8'h3C;
DFS[16'h1662] = 8'h97;
DFS[16'h1663] = 8'hA2;
DFS[16'h1664] = 8'h05;
DFS[16'h1665] = 8'h20;
DFS[16'h1666] = 8'h3C;
DFS[16'h1667] = 8'h97;
DFS[16'h1668] = 8'hD0;
DFS[16'h1669] = 8'hEC;
DFS[16'h166A] = 8'h18;
DFS[16'h166B] = 8'h08;
DFS[16'h166C] = 8'h20;
DFS[16'h166D] = 8'h48;
DFS[16'h166E] = 8'h97;
DFS[16'h166F] = 8'hA2;
DFS[16'h1670] = 8'h05;
DFS[16'h1671] = 8'h20;
DFS[16'h1672] = 8'h3C;
DFS[16'h1673] = 8'h97;
DFS[16'h1674] = 8'hA0;
DFS[16'h1675] = 8'h0C;
DFS[16'h1676] = 8'h20;
DFS[16'h1677] = 8'h56;
DFS[16'h1678] = 8'h97;
DFS[16'h1679] = 8'hB9;
DFS[16'h167A] = 8'h60;
DFS[16'h167B] = 8'h10;
DFS[16'h167C] = 8'h91;
DFS[16'h167D] = 8'hB4;
DFS[16'h167E] = 8'h88;
DFS[16'h167F] = 8'h10;
DFS[16'h1680] = 8'hF8;
DFS[16'h1681] = 8'h28;
DFS[16'h1682] = 8'h60;
DFS[16'h1683] = 8'h20;
DFS[16'h1684] = 8'h4D;
DFS[16'h1685] = 8'h83;
DFS[16'h1686] = 8'h20;
DFS[16'h1687] = 8'h4D;
DFS[16'h1688] = 8'hAB;
DFS[16'h1689] = 8'hA9;
DFS[16'h168A] = 8'h95;
DFS[16'h168B] = 8'h8D;
DFS[16'h168C] = 8'hD8;
DFS[16'h168D] = 8'h10;
DFS[16'h168E] = 8'hA9;
DFS[16'h168F] = 8'h96;
DFS[16'h1690] = 8'h8D;
DFS[16'h1691] = 8'hD9;
DFS[16'h1692] = 8'h10;
DFS[16'h1693] = 8'hD0;
DFS[16'h1694] = 8'hBC;
DFS[16'h1695] = 8'hAC;
DFS[16'h1696] = 8'h69;
DFS[16'h1697] = 8'h10;
DFS[16'h1698] = 8'hCC;
DFS[16'h1699] = 8'h05;
DFS[16'h169A] = 8'h0F;
DFS[16'h169B] = 8'hB0;
DFS[16'h169C] = 8'h28;
DFS[16'h169D] = 8'hB9;
DFS[16'h169E] = 8'h0F;
DFS[16'h169F] = 8'h0E;
DFS[16'h16A0] = 8'h20;
DFS[16'h16A1] = 8'hEE;
DFS[16'h16A2] = 8'h82;
DFS[16'h16A3] = 8'h45;
DFS[16'h16A4] = 8'hCE;
DFS[16'h16A5] = 8'hB0;
DFS[16'h16A6] = 8'h02;
DFS[16'h16A7] = 8'h29;
DFS[16'h16A8] = 8'hDF;
DFS[16'h16A9] = 8'h29;
DFS[16'h16AA] = 8'h7F;
DFS[16'h16AB] = 8'hF0;
DFS[16'h16AC] = 8'h05;
DFS[16'h16AD] = 8'h20;
DFS[16'h16AE] = 8'h10;
DFS[16'h16AF] = 8'h82;
DFS[16'h16B0] = 8'hD0;
DFS[16'h16B1] = 8'hE6;
DFS[16'h16B2] = 8'hA9;
DFS[16'h16B3] = 8'h07;
DFS[16'h16B4] = 8'h20;
DFS[16'h16B5] = 8'h6A;
DFS[16'h16B6] = 8'h97;
DFS[16'h16B7] = 8'h85;
DFS[16'h16B8] = 8'hB0;
DFS[16'h16B9] = 8'hB9;
DFS[16'h16BA] = 8'h08;
DFS[16'h16BB] = 8'h0E;
DFS[16'h16BC] = 8'h20;
DFS[16'h16BD] = 8'h6A;
DFS[16'h16BE] = 8'h97;
DFS[16'h16BF] = 8'hC8;
DFS[16'h16C0] = 8'hC6;
DFS[16'h16C1] = 8'hB0;
DFS[16'h16C2] = 8'hD0;
DFS[16'h16C3] = 8'hF5;
DFS[16'h16C4] = 8'h18;
DFS[16'h16C5] = 8'h8C;
DFS[16'h16C6] = 8'h69;
DFS[16'h16C7] = 8'h10;
DFS[16'h16C8] = 8'hAD;
DFS[16'h16C9] = 8'h04;
DFS[16'h16CA] = 8'h0F;
DFS[16'h16CB] = 8'h8D;
DFS[16'h16CC] = 8'h60;
DFS[16'h16CD] = 8'h10;
DFS[16'h16CE] = 8'h60;
DFS[16'h16CF] = 8'h20;
DFS[16'h16D0] = 8'h4D;
DFS[16'h16D1] = 8'h83;
DFS[16'h16D2] = 8'h20;
DFS[16'h16D3] = 8'h4D;
DFS[16'h16D4] = 8'hAB;
DFS[16'h16D5] = 8'hA9;
DFS[16'h16D6] = 8'h0C;
DFS[16'h16D7] = 8'h20;
DFS[16'h16D8] = 8'h6A;
DFS[16'h16D9] = 8'h97;
DFS[16'h16DA] = 8'hA0;
DFS[16'h16DB] = 8'h00;
DFS[16'h16DC] = 8'hB9;
DFS[16'h16DD] = 8'h00;
DFS[16'h16DE] = 8'h0E;
DFS[16'h16DF] = 8'h20;
DFS[16'h16E0] = 8'h6A;
DFS[16'h16E1] = 8'h97;
DFS[16'h16E2] = 8'hC8;
DFS[16'h16E3] = 8'hC0;
DFS[16'h16E4] = 8'h08;
DFS[16'h16E5] = 8'hD0;
DFS[16'h16E6] = 8'hF5;
DFS[16'h16E7] = 8'hB9;
DFS[16'h16E8] = 8'hF8;
DFS[16'h16E9] = 8'h0E;
DFS[16'h16EA] = 8'h20;
DFS[16'h16EB] = 8'h6A;
DFS[16'h16EC] = 8'h97;
DFS[16'h16ED] = 8'hC8;
DFS[16'h16EE] = 8'hC0;
DFS[16'h16EF] = 8'h0C;
DFS[16'h16F0] = 8'hD0;
DFS[16'h16F1] = 8'hF5;
DFS[16'h16F2] = 8'hAD;
DFS[16'h16F3] = 8'h06;
DFS[16'h16F4] = 8'h0F;
DFS[16'h16F5] = 8'h20;
DFS[16'h16F6] = 8'h05;
DFS[16'h16F7] = 8'h82;
DFS[16'h16F8] = 8'h20;
DFS[16'h16F9] = 8'h6A;
DFS[16'h16FA] = 8'h97;
DFS[16'h16FB] = 8'hA5;
DFS[16'h16FC] = 8'hCF;
DFS[16'h16FD] = 8'h4C;
DFS[16'h16FE] = 8'h6A;
DFS[16'h16FF] = 8'h97;
DFS[16'h1700] = 8'h20;
DFS[16'h1701] = 8'h61;
DFS[16'h1702] = 8'h97;
DFS[16'h1703] = 8'hAD;
DFS[16'h1704] = 8'hCB;
DFS[16'h1705] = 8'h10;
DFS[16'h1706] = 8'h09;
DFS[16'h1707] = 8'h30;
DFS[16'h1708] = 8'h20;
DFS[16'h1709] = 8'h6A;
DFS[16'h170A] = 8'h97;
DFS[16'h170B] = 8'h20;
DFS[16'h170C] = 8'h61;
DFS[16'h170D] = 8'h97;
DFS[16'h170E] = 8'hAD;
DFS[16'h170F] = 8'hCA;
DFS[16'h1710] = 8'h10;
DFS[16'h1711] = 8'h4C;
DFS[16'h1712] = 8'h6A;
DFS[16'h1713] = 8'h97;
DFS[16'h1714] = 8'h20;
DFS[16'h1715] = 8'h61;
DFS[16'h1716] = 8'h97;
DFS[16'h1717] = 8'hAD;
DFS[16'h1718] = 8'hCD;
DFS[16'h1719] = 8'h10;
DFS[16'h171A] = 8'h09;
DFS[16'h171B] = 8'h30;
DFS[16'h171C] = 8'h20;
DFS[16'h171D] = 8'h6A;
DFS[16'h171E] = 8'h97;
DFS[16'h171F] = 8'h20;
DFS[16'h1720] = 8'h61;
DFS[16'h1721] = 8'h97;
DFS[16'h1722] = 8'hAD;
DFS[16'h1723] = 8'hCC;
DFS[16'h1724] = 8'h10;
DFS[16'h1725] = 8'h4C;
DFS[16'h1726] = 8'h6A;
DFS[16'h1727] = 8'h97;
DFS[16'h1728] = 8'h48;
DFS[16'h1729] = 8'hAD;
DFS[16'h172A] = 8'h61;
DFS[16'h172B] = 8'h10;
DFS[16'h172C] = 8'h85;
DFS[16'h172D] = 8'hB8;
DFS[16'h172E] = 8'hAD;
DFS[16'h172F] = 8'h62;
DFS[16'h1730] = 8'h10;
DFS[16'h1731] = 8'h85;
DFS[16'h1732] = 8'hB9;
DFS[16'h1733] = 8'hA2;
DFS[16'h1734] = 8'h00;
DFS[16'h1735] = 8'h68;
DFS[16'h1736] = 8'h60;
DFS[16'h1737] = 8'h20;
DFS[16'h1738] = 8'hE1;
DFS[16'h1739] = 8'h83;
DFS[16'h173A] = 8'hA2;
DFS[16'h173B] = 8'h01;
DFS[16'h173C] = 8'hA0;
DFS[16'h173D] = 8'h04;
DFS[16'h173E] = 8'hFE;
DFS[16'h173F] = 8'h60;
DFS[16'h1740] = 8'h10;
DFS[16'h1741] = 8'hD0;
DFS[16'h1742] = 8'h04;
DFS[16'h1743] = 8'hE8;
DFS[16'h1744] = 8'h88;
DFS[16'h1745] = 8'hD0;
DFS[16'h1746] = 8'hF7;
DFS[16'h1747] = 8'h60;
DFS[16'h1748] = 8'hA2;
DFS[16'h1749] = 8'h03;
DFS[16'h174A] = 8'hA9;
DFS[16'h174B] = 8'hFF;
DFS[16'h174C] = 8'h5D;
DFS[16'h174D] = 8'h65;
DFS[16'h174E] = 8'h10;
DFS[16'h174F] = 8'h9D;
DFS[16'h1750] = 8'h65;
DFS[16'h1751] = 8'h10;
DFS[16'h1752] = 8'hCA;
DFS[16'h1753] = 8'h10;
DFS[16'h1754] = 8'hF5;
DFS[16'h1755] = 8'h60;
DFS[16'h1756] = 8'hAD;
DFS[16'h1757] = 8'h7D;
DFS[16'h1758] = 8'h10;
DFS[16'h1759] = 8'h85;
DFS[16'h175A] = 8'hB4;
DFS[16'h175B] = 8'hAD;
DFS[16'h175C] = 8'h7E;
DFS[16'h175D] = 8'h10;
DFS[16'h175E] = 8'h85;
DFS[16'h175F] = 8'hB5;
DFS[16'h1760] = 8'h60;
DFS[16'h1761] = 8'hA9;
DFS[16'h1762] = 8'h01;
DFS[16'h1763] = 8'hD0;
DFS[16'h1764] = 8'h05;
DFS[16'h1765] = 8'h20;
DFS[16'h1766] = 8'hC1;
DFS[16'h1767] = 8'h90;
DFS[16'h1768] = 8'hB0;
DFS[16'h1769] = 8'hF6;
DFS[16'h176A] = 8'h2C;
DFS[16'h176B] = 8'h81;
DFS[16'h176C] = 8'h10;
DFS[16'h176D] = 8'h10;
DFS[16'h176E] = 8'h06;
DFS[16'h176F] = 8'h8D;
DFS[16'h1770] = 8'hE5;
DFS[16'h1771] = 8'hFE;
DFS[16'h1772] = 8'h4C;
DFS[16'h1773] = 8'h37;
DFS[16'h1774] = 8'h97;
DFS[16'h1775] = 8'h20;
DFS[16'h1776] = 8'h28;
DFS[16'h1777] = 8'h97;
DFS[16'h1778] = 8'h81;
DFS[16'h1779] = 8'hB8;
DFS[16'h177A] = 8'h4C;
DFS[16'h177B] = 8'h37;
DFS[16'h177C] = 8'h97;
DFS[16'h177D] = 8'h20;
DFS[16'h177E] = 8'h85;
DFS[16'h177F] = 8'h97;
DFS[16'h1780] = 8'h20;
DFS[16'h1781] = 8'hAA;
DFS[16'h1782] = 8'h91;
DFS[16'h1783] = 8'h18;
DFS[16'h1784] = 8'h60;
DFS[16'h1785] = 8'h2C;
DFS[16'h1786] = 8'h81;
DFS[16'h1787] = 8'h10;
DFS[16'h1788] = 8'h10;
DFS[16'h1789] = 8'h06;
DFS[16'h178A] = 8'hAD;
DFS[16'h178B] = 8'hE5;
DFS[16'h178C] = 8'hFE;
DFS[16'h178D] = 8'h4C;
DFS[16'h178E] = 8'h37;
DFS[16'h178F] = 8'h97;
DFS[16'h1790] = 8'h20;
DFS[16'h1791] = 8'h28;
DFS[16'h1792] = 8'h97;
DFS[16'h1793] = 8'hA1;
DFS[16'h1794] = 8'hB8;
DFS[16'h1795] = 8'h4C;
DFS[16'h1796] = 8'h37;
DFS[16'h1797] = 8'h97;
DFS[16'h1798] = 8'h2C;
DFS[16'h1799] = 8'hC8;
DFS[16'h179A] = 8'h10;
DFS[16'h179B] = 8'h30;
DFS[16'h179C] = 8'h03;
DFS[16'h179D] = 8'hCE;
DFS[16'h179E] = 8'hC8;
DFS[16'h179F] = 8'h10;
DFS[16'h17A0] = 8'h60;
DFS[16'h17A1] = 8'h20;
DFS[16'h17A2] = 8'h5A;
DFS[16'h17A3] = 8'h98;
DFS[16'h17A4] = 8'h20;
DFS[16'h17A5] = 8'h7E;
DFS[16'h17A6] = 8'h83;
DFS[16'h17A7] = 8'hA9;
DFS[16'h17A8] = 8'h01;
DFS[16'h17A9] = 8'h60;
DFS[16'h17AA] = 8'h20;
DFS[16'h17AB] = 8'h37;
DFS[16'h17AC] = 8'h98;
DFS[16'h17AD] = 8'h20;
DFS[16'h17AE] = 8'h7E;
DFS[16'h17AF] = 8'h83;
DFS[16'h17B0] = 8'h20;
DFS[16'h17B1] = 8'hD1;
DFS[16'h17B2] = 8'h82;
DFS[16'h17B3] = 8'h90;
DFS[16'h17B4] = 8'h24;
DFS[16'h17B5] = 8'h20;
DFS[16'h17B6] = 8'h37;
DFS[16'h17B7] = 8'h98;
DFS[16'h17B8] = 8'h20;
DFS[16'h17B9] = 8'hDF;
DFS[16'h17BA] = 8'h97;
DFS[16'h17BB] = 8'h20;
DFS[16'h17BC] = 8'hFB;
DFS[16'h17BD] = 8'h97;
DFS[16'h17BE] = 8'h50;
DFS[16'h17BF] = 8'h16;
DFS[16'h17C0] = 8'h20;
DFS[16'h17C1] = 8'h37;
DFS[16'h17C2] = 8'h98;
DFS[16'h17C3] = 8'h20;
DFS[16'h17C4] = 8'hDF;
DFS[16'h17C5] = 8'h97;
DFS[16'h17C6] = 8'h50;
DFS[16'h17C7] = 8'h11;
DFS[16'h17C8] = 8'h20;
DFS[16'h17C9] = 8'h37;
DFS[16'h17CA] = 8'h98;
DFS[16'h17CB] = 8'h20;
DFS[16'h17CC] = 8'hFB;
DFS[16'h17CD] = 8'h97;
DFS[16'h17CE] = 8'h50;
DFS[16'h17CF] = 8'h09;
DFS[16'h17D0] = 8'h20;
DFS[16'h17D1] = 8'h5A;
DFS[16'h17D2] = 8'h98;
DFS[16'h17D3] = 8'h20;
DFS[16'h17D4] = 8'h4F;
DFS[16'h17D5] = 8'h98;
DFS[16'h17D6] = 8'h20;
DFS[16'h17D7] = 8'h1E;
DFS[16'h17D8] = 8'h98;
DFS[16'h17D9] = 8'h20;
DFS[16'h17DA] = 8'hC3;
DFS[16'h17DB] = 8'h88;
DFS[16'h17DC] = 8'hA9;
DFS[16'h17DD] = 8'h01;
DFS[16'h17DE] = 8'h60;
DFS[16'h17DF] = 8'h20;
DFS[16'h17E0] = 8'hE1;
DFS[16'h17E1] = 8'h83;
DFS[16'h17E2] = 8'hA0;
DFS[16'h17E3] = 8'h02;
DFS[16'h17E4] = 8'hB1;
DFS[16'h17E5] = 8'hB0;
DFS[16'h17E6] = 8'h9D;
DFS[16'h17E7] = 8'h08;
DFS[16'h17E8] = 8'h0F;
DFS[16'h17E9] = 8'hC8;
DFS[16'h17EA] = 8'hB1;
DFS[16'h17EB] = 8'hB0;
DFS[16'h17EC] = 8'h9D;
DFS[16'h17ED] = 8'h09;
DFS[16'h17EE] = 8'h0F;
DFS[16'h17EF] = 8'hC8;
DFS[16'h17F0] = 8'hB1;
DFS[16'h17F1] = 8'hB0;
DFS[16'h17F2] = 8'h0A;
DFS[16'h17F3] = 8'h0A;
DFS[16'h17F4] = 8'h5D;
DFS[16'h17F5] = 8'h0E;
DFS[16'h17F6] = 8'h0F;
DFS[16'h17F7] = 8'h29;
DFS[16'h17F8] = 8'h0C;
DFS[16'h17F9] = 8'h10;
DFS[16'h17FA] = 8'h1B;
DFS[16'h17FB] = 8'h20;
DFS[16'h17FC] = 8'hE1;
DFS[16'h17FD] = 8'h83;
DFS[16'h17FE] = 8'hA0;
DFS[16'h17FF] = 8'h06;
DFS[16'h1800] = 8'hB1;
DFS[16'h1801] = 8'hB0;
DFS[16'h1802] = 8'h9D;
DFS[16'h1803] = 8'h0A;
DFS[16'h1804] = 8'h0F;
DFS[16'h1805] = 8'hC8;
DFS[16'h1806] = 8'hB1;
DFS[16'h1807] = 8'hB0;
DFS[16'h1808] = 8'h9D;
DFS[16'h1809] = 8'h0B;
DFS[16'h180A] = 8'h0F;
DFS[16'h180B] = 8'hC8;
DFS[16'h180C] = 8'hB1;
DFS[16'h180D] = 8'hB0;
DFS[16'h180E] = 8'h6A;
DFS[16'h180F] = 8'h6A;
DFS[16'h1810] = 8'h6A;
DFS[16'h1811] = 8'h5D;
DFS[16'h1812] = 8'h0E;
DFS[16'h1813] = 8'h0F;
DFS[16'h1814] = 8'h29;
DFS[16'h1815] = 8'hC0;
DFS[16'h1816] = 8'h5D;
DFS[16'h1817] = 8'h0E;
DFS[16'h1818] = 8'h0F;
DFS[16'h1819] = 8'h9D;
DFS[16'h181A] = 8'h0E;
DFS[16'h181B] = 8'h0F;
DFS[16'h181C] = 8'hB8;
DFS[16'h181D] = 8'h60;
DFS[16'h181E] = 8'h20;
DFS[16'h181F] = 8'hE1;
DFS[16'h1820] = 8'h83;
DFS[16'h1821] = 8'hA0;
DFS[16'h1822] = 8'h0E;
DFS[16'h1823] = 8'hB1;
DFS[16'h1824] = 8'hB0;
DFS[16'h1825] = 8'h29;
DFS[16'h1826] = 8'h0A;
DFS[16'h1827] = 8'hF0;
DFS[16'h1828] = 8'h02;
DFS[16'h1829] = 8'hA9;
DFS[16'h182A] = 8'h80;
DFS[16'h182B] = 8'h5D;
DFS[16'h182C] = 8'h0F;
DFS[16'h182D] = 8'h0E;
DFS[16'h182E] = 8'h29;
DFS[16'h182F] = 8'h80;
DFS[16'h1830] = 8'h5D;
DFS[16'h1831] = 8'h0F;
DFS[16'h1832] = 8'h0E;
DFS[16'h1833] = 8'h9D;
DFS[16'h1834] = 8'h0F;
DFS[16'h1835] = 8'h0E;
DFS[16'h1836] = 8'h60;
DFS[16'h1837] = 8'h20;
DFS[16'h1838] = 8'h64;
DFS[16'h1839] = 8'h98;
DFS[16'h183A] = 8'h90;
DFS[16'h183B] = 8'h23;
DFS[16'h183C] = 8'hB9;
DFS[16'h183D] = 8'h0F;
DFS[16'h183E] = 8'h0E;
DFS[16'h183F] = 8'h10;
DFS[16'h1840] = 8'h22;
DFS[16'h1841] = 8'h20;
DFS[16'h1842] = 8'h2B;
DFS[16'h1843] = 8'h80;
DFS[16'h1844] = 8'hC3;
DFS[16'h1845] = 8'h6C;
DFS[16'h1846] = 8'h6F;
DFS[16'h1847] = 8'h63;
DFS[16'h1848] = 8'h6B;
DFS[16'h1849] = 8'h65;
DFS[16'h184A] = 8'h64;
DFS[16'h184B] = 8'h00;
DFS[16'h184C] = 8'h20;
DFS[16'h184D] = 8'h3C;
DFS[16'h184E] = 8'h98;
DFS[16'h184F] = 8'h20;
DFS[16'h1850] = 8'hE1;
DFS[16'h1851] = 8'h83;
DFS[16'h1852] = 8'h20;
DFS[16'h1853] = 8'h9E;
DFS[16'h1854] = 8'h8F;
DFS[16'h1855] = 8'h90;
DFS[16'h1856] = 8'h21;
DFS[16'h1857] = 8'h4C;
DFS[16'h1858] = 8'h02;
DFS[16'h1859] = 8'h8F;
DFS[16'h185A] = 8'h20;
DFS[16'h185B] = 8'h64;
DFS[16'h185C] = 8'h98;
DFS[16'h185D] = 8'hB0;
DFS[16'h185E] = 8'h19;
DFS[16'h185F] = 8'h68;
DFS[16'h1860] = 8'h68;
DFS[16'h1861] = 8'hA9;
DFS[16'h1862] = 8'h00;
DFS[16'h1863] = 8'h60;
DFS[16'h1864] = 8'h20;
DFS[16'h1865] = 8'h06;
DFS[16'h1866] = 8'h81;
DFS[16'h1867] = 8'h20;
DFS[16'h1868] = 8'h96;
DFS[16'h1869] = 8'h82;
DFS[16'h186A] = 8'h90;
DFS[16'h186B] = 8'h0C;
DFS[16'h186C] = 8'h98;
DFS[16'h186D] = 8'hAA;
DFS[16'h186E] = 8'hAD;
DFS[16'h186F] = 8'hDC;
DFS[16'h1870] = 8'h10;
DFS[16'h1871] = 8'h85;
DFS[16'h1872] = 8'hB0;
DFS[16'h1873] = 8'hAD;
DFS[16'h1874] = 8'hDD;
DFS[16'h1875] = 8'h10;
DFS[16'h1876] = 8'h85;
DFS[16'h1877] = 8'hB1;
DFS[16'h1878] = 8'h60;
DFS[16'h1879] = 8'hA9;
DFS[16'h187A] = 8'h83;
DFS[16'h187B] = 8'h20;
DFS[16'h187C] = 8'hF4;
DFS[16'h187D] = 8'hFF;
DFS[16'h187E] = 8'h8C;
DFS[16'h187F] = 8'hD0;
DFS[16'h1880] = 8'h10;
DFS[16'h1881] = 8'hA9;
DFS[16'h1882] = 8'h84;
DFS[16'h1883] = 8'h20;
DFS[16'h1884] = 8'hF4;
DFS[16'h1885] = 8'hFF;
DFS[16'h1886] = 8'h98;
DFS[16'h1887] = 8'h38;
DFS[16'h1888] = 8'hED;
DFS[16'h1889] = 8'hD0;
DFS[16'h188A] = 8'h10;
DFS[16'h188B] = 8'h8D;
DFS[16'h188C] = 8'hD1;
DFS[16'h188D] = 8'h10;
DFS[16'h188E] = 8'h60;
DFS[16'h188F] = 8'hA2;
DFS[16'h1890] = 8'h0A;
DFS[16'h1891] = 8'h20;
DFS[16'h1892] = 8'h2C;
DFS[16'h1893] = 8'h99;
DFS[16'h1894] = 8'h20;
DFS[16'h1895] = 8'h9E;
DFS[16'h1896] = 8'h98;
DFS[16'h1897] = 8'hA0;
DFS[16'h1898] = 8'hD5;
DFS[16'h1899] = 8'hA9;
DFS[16'h189A] = 8'hFF;
DFS[16'h189B] = 8'h91;
DFS[16'h189C] = 8'hB0;
DFS[16'h189D] = 8'h60;
DFS[16'h189E] = 8'h48;
DFS[16'h189F] = 8'hA6;
DFS[16'h18A0] = 8'hF4;
DFS[16'h18A1] = 8'hA9;
DFS[16'h18A2] = 8'h00;
DFS[16'h18A3] = 8'h85;
DFS[16'h18A4] = 8'hB0;
DFS[16'h18A5] = 8'hBD;
DFS[16'h18A6] = 8'hF0;
DFS[16'h18A7] = 8'h0D;
DFS[16'h18A8] = 8'h85;
DFS[16'h18A9] = 8'hB1;
DFS[16'h18AA] = 8'h68;
DFS[16'h18AB] = 8'h60;
DFS[16'h18AC] = 8'h00;
DFS[16'h18AD] = 8'h00;
DFS[16'h18AE] = 8'h00;
DFS[16'h18AF] = 8'h00;
DFS[16'h18B0] = 8'h00;
DFS[16'h18B1] = 8'h00;
DFS[16'h18B2] = 8'h00;
DFS[16'h18B3] = 8'h00;
DFS[16'h18B4] = 8'h00;
DFS[16'h18B5] = 8'h00;
DFS[16'h18B6] = 8'h00;
DFS[16'h18B7] = 8'h00;
DFS[16'h18B8] = 8'h00;
DFS[16'h18B9] = 8'h00;
DFS[16'h18BA] = 8'h00;
DFS[16'h18BB] = 8'h00;
DFS[16'h18BC] = 8'h00;
DFS[16'h18BD] = 8'h00;
DFS[16'h18BE] = 8'h00;
DFS[16'h18BF] = 8'h00;
DFS[16'h18C0] = 8'h00;
DFS[16'h18C1] = 8'h00;
DFS[16'h18C2] = 8'h00;
DFS[16'h18C3] = 8'h00;
DFS[16'h18C4] = 8'h00;
DFS[16'h18C5] = 8'h00;
DFS[16'h18C6] = 8'h00;
DFS[16'h18C7] = 8'h00;
DFS[16'h18C8] = 8'h00;
DFS[16'h18C9] = 8'h00;
DFS[16'h18CA] = 8'h00;
DFS[16'h18CB] = 8'h00;
DFS[16'h18CC] = 8'h00;
DFS[16'h18CD] = 8'h00;
DFS[16'h18CE] = 8'h00;
DFS[16'h18CF] = 8'h00;
DFS[16'h18D0] = 8'h00;
DFS[16'h18D1] = 8'h00;
DFS[16'h18D2] = 8'h00;
DFS[16'h18D3] = 8'h00;
DFS[16'h18D4] = 8'h00;
DFS[16'h18D5] = 8'h00;
DFS[16'h18D6] = 8'h00;
DFS[16'h18D7] = 8'h00;
DFS[16'h18D8] = 8'h00;
DFS[16'h18D9] = 8'h00;
DFS[16'h18DA] = 8'h00;
DFS[16'h18DB] = 8'h00;
DFS[16'h18DC] = 8'h00;
DFS[16'h18DD] = 8'h00;
DFS[16'h18DE] = 8'h00;
DFS[16'h18DF] = 8'h00;
DFS[16'h18E0] = 8'h00;
DFS[16'h18E1] = 8'h00;
DFS[16'h18E2] = 8'h00;
DFS[16'h18E3] = 8'h00;
DFS[16'h18E4] = 8'h00;
DFS[16'h18E5] = 8'h00;
DFS[16'h18E6] = 8'h00;
DFS[16'h18E7] = 8'h00;
DFS[16'h18E8] = 8'h00;
DFS[16'h18E9] = 8'h00;
DFS[16'h18EA] = 8'h00;
DFS[16'h18EB] = 8'h00;
DFS[16'h18EC] = 8'h00;
DFS[16'h18ED] = 8'h00;
DFS[16'h18EE] = 8'h00;
DFS[16'h18EF] = 8'h00;
DFS[16'h18F0] = 8'h00;
DFS[16'h18F1] = 8'h00;
DFS[16'h18F2] = 8'h00;
DFS[16'h18F3] = 8'h00;
DFS[16'h18F4] = 8'h00;
DFS[16'h18F5] = 8'h00;
DFS[16'h18F6] = 8'h00;
DFS[16'h18F7] = 8'h00;
DFS[16'h18F8] = 8'h00;
DFS[16'h18F9] = 8'h00;
DFS[16'h18FA] = 8'h00;
DFS[16'h18FB] = 8'h00;
DFS[16'h18FC] = 8'h00;
DFS[16'h18FD] = 8'h00;
DFS[16'h18FE] = 8'h00;
DFS[16'h18FF] = 8'h00;
DFS[16'h1900] = 8'h00;
DFS[16'h1901] = 8'h00;
DFS[16'h1902] = 8'h00;
DFS[16'h1903] = 8'h00;
DFS[16'h1904] = 8'h00;
DFS[16'h1905] = 8'h60;
DFS[16'h1906] = 8'h20;
DFS[16'h1907] = 8'hE1;
DFS[16'h1908] = 8'h83;
DFS[16'h1909] = 8'hA9;
DFS[16'h190A] = 8'h0F;
DFS[16'h190B] = 8'hA2;
DFS[16'h190C] = 8'h01;
DFS[16'h190D] = 8'hA0;
DFS[16'h190E] = 8'h00;
DFS[16'h190F] = 8'hF0;
DFS[16'h1910] = 8'h25;
DFS[16'h1911] = 8'hA9;
DFS[16'h1912] = 8'hC7;
DFS[16'h1913] = 8'hA2;
DFS[16'h1914] = 8'h00;
DFS[16'h1915] = 8'hF0;
DFS[16'h1916] = 8'hF6;
DFS[16'h1917] = 8'hAA;
DFS[16'h1918] = 8'hA9;
DFS[16'h1919] = 8'h03;
DFS[16'h191A] = 8'hD0;
DFS[16'h191B] = 8'h1A;
DFS[16'h191C] = 8'hA9;
DFS[16'h191D] = 8'hEC;
DFS[16'h191E] = 8'hD0;
DFS[16'h191F] = 8'h12;
DFS[16'h1920] = 8'hA9;
DFS[16'h1921] = 8'hC7;
DFS[16'h1922] = 8'hD0;
DFS[16'h1923] = 8'h0E;
DFS[16'h1924] = 8'hA9;
DFS[16'h1925] = 8'hEA;
DFS[16'h1926] = 8'hD0;
DFS[16'h1927] = 8'h0A;
DFS[16'h1928] = 8'hA9;
DFS[16'h1929] = 8'hA8;
DFS[16'h192A] = 8'hD0;
DFS[16'h192B] = 8'h06;
DFS[16'h192C] = 8'hA9;
DFS[16'h192D] = 8'h8F;
DFS[16'h192E] = 8'hD0;
DFS[16'h192F] = 8'h06;
DFS[16'h1930] = 8'hA9;
DFS[16'h1931] = 8'hFF;
DFS[16'h1932] = 8'hA2;
DFS[16'h1933] = 8'h00;
DFS[16'h1934] = 8'hA0;
DFS[16'h1935] = 8'hFF;
DFS[16'h1936] = 8'h4C;
DFS[16'h1937] = 8'hF4;
DFS[16'h1938] = 8'hFF;
DFS[16'h1939] = 8'h4C;
DFS[16'h193A] = 8'h2E;
DFS[16'h193B] = 8'h21;
DFS[16'h193C] = 8'h42;
DFS[16'h193D] = 8'h4F;
DFS[16'h193E] = 8'h4F;
DFS[16'h193F] = 8'h54;
DFS[16'h1940] = 8'h0D;
DFS[16'h1941] = 8'h45;
DFS[16'h1942] = 8'h2E;
DFS[16'h1943] = 8'h21;
DFS[16'h1944] = 8'h42;
DFS[16'h1945] = 8'h4F;
DFS[16'h1946] = 8'h4F;
DFS[16'h1947] = 8'h54;
DFS[16'h1948] = 8'h0D;
DFS[16'h1949] = 8'h1B;
DFS[16'h194A] = 8'hFF;
DFS[16'h194B] = 8'h1E;
DFS[16'h194C] = 8'hFF;
DFS[16'h194D] = 8'h21;
DFS[16'h194E] = 8'hFF;
DFS[16'h194F] = 8'h24;
DFS[16'h1950] = 8'hFF;
DFS[16'h1951] = 8'h27;
DFS[16'h1952] = 8'hFF;
DFS[16'h1953] = 8'h2A;
DFS[16'h1954] = 8'hFF;
DFS[16'h1955] = 8'h2D;
DFS[16'h1956] = 8'hFF;
DFS[16'h1957] = 8'h7B;
DFS[16'h1958] = 8'h95;
DFS[16'h1959] = 8'h00;
DFS[16'h195A] = 8'h07;
DFS[16'h195B] = 8'h90;
DFS[16'h195C] = 8'h00;
DFS[16'h195D] = 8'hC1;
DFS[16'h195E] = 8'h90;
DFS[16'h195F] = 8'h00;
DFS[16'h1960] = 8'hAA;
DFS[16'h1961] = 8'h91;
DFS[16'h1962] = 8'h00;
DFS[16'h1963] = 8'hD0;
DFS[16'h1964] = 8'h95;
DFS[16'h1965] = 8'h00;
DFS[16'h1966] = 8'h93;
DFS[16'h1967] = 8'h8E;
DFS[16'h1968] = 8'h00;
DFS[16'h1969] = 8'hAA;
DFS[16'h196A] = 8'h95;
DFS[16'h196B] = 8'h00;
DFS[16'h196C] = 8'h1B;
DFS[16'h196D] = 8'h8C;
DFS[16'h196E] = 8'hD3;
DFS[16'h196F] = 8'h6B;
DFS[16'h1970] = 8'hD3;
DFS[16'h1971] = 8'h1D;
DFS[16'h1972] = 8'hE1;
DFS[16'h1973] = 8'hDC;
DFS[16'h1974] = 8'h97;
DFS[16'h1975] = 8'h89;
DFS[16'h1976] = 8'h90;
DFS[16'h1977] = 8'h87;
DFS[16'h1978] = 8'h86;
DFS[16'h1979] = 8'h87;
DFS[16'h197A] = 8'h84;
DFS[16'h197B] = 8'h8D;
DFS[16'h197C] = 8'h8D;
DFS[16'h197D] = 8'h97;
DFS[16'h197E] = 8'hF1;
DFS[16'h197F] = 8'h3C;
DFS[16'h1980] = 8'hBC;
DFS[16'h1981] = 8'h8F;
DFS[16'h1982] = 8'h9B;
DFS[16'h1983] = 8'h95;
DFS[16'h1984] = 8'h93;
DFS[16'h1985] = 8'h85;
DFS[16'h1986] = 8'hB4;
DFS[16'h1987] = 8'hBF;
DFS[16'h1988] = 8'hC7;
DFS[16'h1989] = 8'hCF;
DFS[16'h198A] = 8'hA0;
DFS[16'h198B] = 8'hA9;
DFS[16'h198C] = 8'h87;
DFS[16'h198D] = 8'h87;
DFS[16'h198E] = 8'h97;
DFS[16'h198F] = 8'h97;
DFS[16'h1990] = 8'h97;
DFS[16'h1991] = 8'h97;
DFS[16'h1992] = 8'h97;
DFS[16'h1993] = 8'h97;
DFS[16'h1994] = 8'h12;
DFS[16'h1995] = 8'h32;
DFS[16'h1996] = 8'h5D;
DFS[16'h1997] = 8'hCD;
DFS[16'h1998] = 8'hA2;
DFS[16'h1999] = 8'hBD;
DFS[16'h199A] = 8'h87;
DFS[16'h199B] = 8'h8D;
DFS[16'h199C] = 8'h8D;
DFS[16'h199D] = 8'h8D;
DFS[16'h199E] = 8'h8D;
DFS[16'h199F] = 8'h8D;
DFS[16'h19A0] = 8'h8D;
DFS[16'h19A1] = 8'h8D;
DFS[16'h19A2] = 8'h74;
DFS[16'h19A3] = 8'h54;
DFS[16'h19A4] = 8'h00;
DFS[16'h19A5] = 8'h0F;
DFS[16'h19A6] = 8'h1A;
DFS[16'h19A7] = 8'h0F;
DFS[16'h19A8] = 8'h1A;
DFS[16'h19A9] = 8'h63;
DFS[16'h19AA] = 8'h43;
DFS[16'h19AB] = 8'hB7;
DFS[16'h19AC] = 8'h7D;
DFS[16'h19AD] = 8'h7D;
DFS[16'h19AE] = 8'h65;
DFS[16'h19AF] = 8'h65;
DFS[16'h19B0] = 8'hCF;
DFS[16'h19B1] = 8'h00;
DFS[16'h19B2] = 8'h14;
DFS[16'h19B3] = 8'h83;
DFS[16'h19B4] = 8'h85;
DFS[16'h19B5] = 8'h97;
DFS[16'h19B6] = 8'h97;
DFS[16'h19B7] = 8'h97;
DFS[16'h19B8] = 8'h97;
DFS[16'h19B9] = 8'h96;
DFS[16'h19BA] = 8'h97;
DFS[16'h19BB] = 8'h97;
DFS[16'h19BC] = 8'h96;
DFS[16'h19BD] = 8'h04;
DFS[16'h19BE] = 8'h02;
DFS[16'h19BF] = 8'h03;
DFS[16'h19C0] = 8'h06;
DFS[16'h19C1] = 8'h07;
DFS[16'h19C2] = 8'h04;
DFS[16'h19C3] = 8'h04;
DFS[16'h19C4] = 8'h04;
DFS[16'h19C5] = 8'h04;
DFS[16'h19C6] = 8'h98;
DFS[16'h19C7] = 8'hA2;
DFS[16'h19C8] = 8'hFF;
DFS[16'h19C9] = 8'hA0;
DFS[16'h19CA] = 8'h0E;
DFS[16'h19CB] = 8'h48;
DFS[16'h19CC] = 8'h20;
DFS[16'h19CD] = 8'h65;
DFS[16'h19CE] = 8'h80;
DFS[16'h19CF] = 8'h0D;
DFS[16'h19D0] = 8'h44;
DFS[16'h19D1] = 8'h46;
DFS[16'h19D2] = 8'h53;
DFS[16'h19D3] = 8'h20;
DFS[16'h19D4] = 8'h30;
DFS[16'h19D5] = 8'h2E;
DFS[16'h19D6] = 8'h39;
DFS[16'h19D7] = 8'h30;
DFS[16'h19D8] = 8'h0D;
DFS[16'h19D9] = 8'h86;
DFS[16'h19DA] = 8'hB8;
DFS[16'h19DB] = 8'h20;
DFS[16'h19DC] = 8'hCB;
DFS[16'h19DD] = 8'h9F;
DFS[16'h19DE] = 8'h20;
DFS[16'h19DF] = 8'h19;
DFS[16'h19E0] = 8'h9A;
DFS[16'h19E1] = 8'h20;
DFS[16'h19E2] = 8'h9A;
DFS[16'h19E3] = 8'h9F;
DFS[16'h19E4] = 8'h88;
DFS[16'h19E5] = 8'hD0;
DFS[16'h19E6] = 8'hF4;
DFS[16'h19E7] = 8'h68;
DFS[16'h19E8] = 8'hA8;
DFS[16'h19E9] = 8'hA2;
DFS[16'h19EA] = 8'hA0;
DFS[16'h19EB] = 8'h4C;
DFS[16'h19EC] = 8'h71;
DFS[16'h19ED] = 8'h86;
DFS[16'h19EE] = 8'h98;
DFS[16'h19EF] = 8'hA2;
DFS[16'h19F0] = 8'h74;
DFS[16'h19F1] = 8'hA0;
DFS[16'h19F2] = 8'h05;
DFS[16'h19F3] = 8'hD0;
DFS[16'h19F4] = 8'hD6;
DFS[16'h19F5] = 8'h20;
DFS[16'h19F6] = 8'hBF;
DFS[16'h19F7] = 8'h86;
DFS[16'h19F8] = 8'hF0;
DFS[16'h19F9] = 8'h60;
DFS[16'h19FA] = 8'h20;
DFS[16'h19FB] = 8'hC5;
DFS[16'h19FC] = 8'hFF;
DFS[16'h19FD] = 8'h90;
DFS[16'h19FE] = 8'hFB;
DFS[16'h19FF] = 8'hB0;
DFS[16'h1A00] = 8'hE8;
DFS[16'h1A01] = 8'h20;
DFS[16'h1A02] = 8'hBF;
DFS[16'h1A03] = 8'h86;
DFS[16'h1A04] = 8'hD0;
DFS[16'h1A05] = 8'h54;
DFS[16'h1A06] = 8'h20;
DFS[16'h1A07] = 8'h33;
DFS[16'h1A08] = 8'h80;
DFS[16'h1A09] = 8'hDC;
DFS[16'h1A0A] = 8'h53;
DFS[16'h1A0B] = 8'h79;
DFS[16'h1A0C] = 8'h6E;
DFS[16'h1A0D] = 8'h74;
DFS[16'h1A0E] = 8'h61;
DFS[16'h1A0F] = 8'h78;
DFS[16'h1A10] = 8'h3A;
DFS[16'h1A11] = 8'h20;
DFS[16'h1A12] = 8'hEA;
DFS[16'h1A13] = 8'h20;
DFS[16'h1A14] = 8'h19;
DFS[16'h1A15] = 8'h9A;
DFS[16'h1A16] = 8'h4C;
DFS[16'h1A17] = 8'h8A;
DFS[16'h1A18] = 8'h80;
DFS[16'h1A19] = 8'hA6;
DFS[16'h1A1A] = 8'hB8;
DFS[16'h1A1B] = 8'hE8;
DFS[16'h1A1C] = 8'hBD;
DFS[16'h1A1D] = 8'hB8;
DFS[16'h1A1E] = 8'h85;
DFS[16'h1A1F] = 8'h30;
DFS[16'h1A20] = 8'h06;
DFS[16'h1A21] = 8'h20;
DFS[16'h1A22] = 8'h9C;
DFS[16'h1A23] = 8'h80;
DFS[16'h1A24] = 8'h4C;
DFS[16'h1A25] = 8'h1B;
DFS[16'h1A26] = 8'h9A;
DFS[16'h1A27] = 8'hE8;
DFS[16'h1A28] = 8'hE8;
DFS[16'h1A29] = 8'h86;
DFS[16'h1A2A] = 8'hB8;
DFS[16'h1A2B] = 8'hBD;
DFS[16'h1A2C] = 8'hB8;
DFS[16'h1A2D] = 8'h85;
DFS[16'h1A2E] = 8'h20;
DFS[16'h1A2F] = 8'h34;
DFS[16'h1A30] = 8'h9A;
DFS[16'h1A31] = 8'h20;
DFS[16'h1A32] = 8'h05;
DFS[16'h1A33] = 8'h82;
DFS[16'h1A34] = 8'h20;
DFS[16'h1A35] = 8'hE1;
DFS[16'h1A36] = 8'h83;
DFS[16'h1A37] = 8'h29;
DFS[16'h1A38] = 8'h0F;
DFS[16'h1A39] = 8'hF0;
DFS[16'h1A3A] = 8'h1F;
DFS[16'h1A3B] = 8'hA8;
DFS[16'h1A3C] = 8'hA9;
DFS[16'h1A3D] = 8'h20;
DFS[16'h1A3E] = 8'h20;
DFS[16'h1A3F] = 8'h9C;
DFS[16'h1A40] = 8'h80;
DFS[16'h1A41] = 8'hA2;
DFS[16'h1A42] = 8'h00;
DFS[16'h1A43] = 8'hBD;
DFS[16'h1A44] = 8'h5B;
DFS[16'h1A45] = 8'h9A;
DFS[16'h1A46] = 8'hF0;
DFS[16'h1A47] = 8'h03;
DFS[16'h1A48] = 8'hE8;
DFS[16'h1A49] = 8'hD0;
DFS[16'h1A4A] = 8'hF8;
DFS[16'h1A4B] = 8'h88;
DFS[16'h1A4C] = 8'hD0;
DFS[16'h1A4D] = 8'hFA;
DFS[16'h1A4E] = 8'hE8;
DFS[16'h1A4F] = 8'hBD;
DFS[16'h1A50] = 8'h5B;
DFS[16'h1A51] = 8'h9A;
DFS[16'h1A52] = 8'hF0;
DFS[16'h1A53] = 8'h06;
DFS[16'h1A54] = 8'h20;
DFS[16'h1A55] = 8'h9C;
DFS[16'h1A56] = 8'h80;
DFS[16'h1A57] = 8'h4C;
DFS[16'h1A58] = 8'h4E;
DFS[16'h1A59] = 8'h9A;
DFS[16'h1A5A] = 8'h60;
DFS[16'h1A5B] = 8'h00;
DFS[16'h1A5C] = 8'h3C;
DFS[16'h1A5D] = 8'h66;
DFS[16'h1A5E] = 8'h73;
DFS[16'h1A5F] = 8'h70;
DFS[16'h1A60] = 8'h3E;
DFS[16'h1A61] = 8'h00;
DFS[16'h1A62] = 8'h3C;
DFS[16'h1A63] = 8'h61;
DFS[16'h1A64] = 8'h66;
DFS[16'h1A65] = 8'h73;
DFS[16'h1A66] = 8'h70;
DFS[16'h1A67] = 8'h3E;
DFS[16'h1A68] = 8'h00;
DFS[16'h1A69] = 8'h28;
DFS[16'h1A6A] = 8'h4C;
DFS[16'h1A6B] = 8'h29;
DFS[16'h1A6C] = 8'h00;
DFS[16'h1A6D] = 8'h3C;
DFS[16'h1A6E] = 8'h73;
DFS[16'h1A6F] = 8'h72;
DFS[16'h1A70] = 8'h63;
DFS[16'h1A71] = 8'h20;
DFS[16'h1A72] = 8'h64;
DFS[16'h1A73] = 8'h72;
DFS[16'h1A74] = 8'h76;
DFS[16'h1A75] = 8'h3E;
DFS[16'h1A76] = 8'h00;
DFS[16'h1A77] = 8'h3C;
DFS[16'h1A78] = 8'h64;
DFS[16'h1A79] = 8'h65;
DFS[16'h1A7A] = 8'h73;
DFS[16'h1A7B] = 8'h74;
DFS[16'h1A7C] = 8'h20;
DFS[16'h1A7D] = 8'h64;
DFS[16'h1A7E] = 8'h72;
DFS[16'h1A7F] = 8'h76;
DFS[16'h1A80] = 8'h3E;
DFS[16'h1A81] = 8'h00;
DFS[16'h1A82] = 8'h3C;
DFS[16'h1A83] = 8'h64;
DFS[16'h1A84] = 8'h65;
DFS[16'h1A85] = 8'h73;
DFS[16'h1A86] = 8'h74;
DFS[16'h1A87] = 8'h20;
DFS[16'h1A88] = 8'h64;
DFS[16'h1A89] = 8'h72;
DFS[16'h1A8A] = 8'h76;
DFS[16'h1A8B] = 8'h3E;
DFS[16'h1A8C] = 8'h20;
DFS[16'h1A8D] = 8'h3C;
DFS[16'h1A8E] = 8'h61;
DFS[16'h1A8F] = 8'h66;
DFS[16'h1A90] = 8'h73;
DFS[16'h1A91] = 8'h70;
DFS[16'h1A92] = 8'h3E;
DFS[16'h1A93] = 8'h00;
DFS[16'h1A94] = 8'h3C;
DFS[16'h1A95] = 8'h6F;
DFS[16'h1A96] = 8'h6C;
DFS[16'h1A97] = 8'h64;
DFS[16'h1A98] = 8'h20;
DFS[16'h1A99] = 8'h66;
DFS[16'h1A9A] = 8'h73;
DFS[16'h1A9B] = 8'h70;
DFS[16'h1A9C] = 8'h3E;
DFS[16'h1A9D] = 8'h00;
DFS[16'h1A9E] = 8'h3C;
DFS[16'h1A9F] = 8'h6E;
DFS[16'h1AA0] = 8'h65;
DFS[16'h1AA1] = 8'h77;
DFS[16'h1AA2] = 8'h20;
DFS[16'h1AA3] = 8'h66;
DFS[16'h1AA4] = 8'h73;
DFS[16'h1AA5] = 8'h70;
DFS[16'h1AA6] = 8'h3E;
DFS[16'h1AA7] = 8'h00;
DFS[16'h1AA8] = 8'h28;
DFS[16'h1AA9] = 8'h3C;
DFS[16'h1AAA] = 8'h64;
DFS[16'h1AAB] = 8'h69;
DFS[16'h1AAC] = 8'h72;
DFS[16'h1AAD] = 8'h3E;
DFS[16'h1AAE] = 8'h29;
DFS[16'h1AAF] = 8'h00;
DFS[16'h1AB0] = 8'h28;
DFS[16'h1AB1] = 8'h3C;
DFS[16'h1AB2] = 8'h64;
DFS[16'h1AB3] = 8'h72;
DFS[16'h1AB4] = 8'h76;
DFS[16'h1AB5] = 8'h3E;
DFS[16'h1AB6] = 8'h29;
DFS[16'h1AB7] = 8'h00;
DFS[16'h1AB8] = 8'h3C;
DFS[16'h1AB9] = 8'h74;
DFS[16'h1ABA] = 8'h69;
DFS[16'h1ABB] = 8'h74;
DFS[16'h1ABC] = 8'h6C;
DFS[16'h1ABD] = 8'h65;
DFS[16'h1ABE] = 8'h3E;
DFS[16'h1ABF] = 8'h00;
DFS[16'h1AC0] = 8'h20;
DFS[16'h1AC1] = 8'h58;
DFS[16'h1AC2] = 8'h83;
DFS[16'h1AC3] = 8'h20;
DFS[16'h1AC4] = 8'h65;
DFS[16'h1AC5] = 8'h80;
DFS[16'h1AC6] = 8'h43;
DFS[16'h1AC7] = 8'h6F;
DFS[16'h1AC8] = 8'h6D;
DFS[16'h1AC9] = 8'h70;
DFS[16'h1ACA] = 8'h61;
DFS[16'h1ACB] = 8'h63;
DFS[16'h1ACC] = 8'h74;
DFS[16'h1ACD] = 8'h69;
DFS[16'h1ACE] = 8'h6E;
DFS[16'h1ACF] = 8'h67;
DFS[16'h1AD0] = 8'h20;
DFS[16'h1AD1] = 8'h64;
DFS[16'h1AD2] = 8'h72;
DFS[16'h1AD3] = 8'h69;
DFS[16'h1AD4] = 8'h76;
DFS[16'h1AD5] = 8'h65;
DFS[16'h1AD6] = 8'h20;
DFS[16'h1AD7] = 8'h8D;
DFS[16'h1AD8] = 8'hD2;
DFS[16'h1AD9] = 8'h10;
DFS[16'h1ADA] = 8'h8D;
DFS[16'h1ADB] = 8'hD3;
DFS[16'h1ADC] = 8'h10;
DFS[16'h1ADD] = 8'h20;
DFS[16'h1ADE] = 8'hCA;
DFS[16'h1ADF] = 8'h80;
DFS[16'h1AE0] = 8'h20;
DFS[16'h1AE1] = 8'h9A;
DFS[16'h1AE2] = 8'h9F;
DFS[16'h1AE3] = 8'hA0;
DFS[16'h1AE4] = 8'h00;
DFS[16'h1AE5] = 8'h20;
DFS[16'h1AE6] = 8'h05;
DFS[16'h1AE7] = 8'h8E;
DFS[16'h1AE8] = 8'h20;
DFS[16'h1AE9] = 8'h79;
DFS[16'h1AEA] = 8'h98;
DFS[16'h1AEB] = 8'h20;
DFS[16'h1AEC] = 8'h47;
DFS[16'h1AED] = 8'h83;
DFS[16'h1AEE] = 8'hAC;
DFS[16'h1AEF] = 8'h05;
DFS[16'h1AF0] = 8'h0F;
DFS[16'h1AF1] = 8'h84;
DFS[16'h1AF2] = 8'hCC;
DFS[16'h1AF3] = 8'hA9;
DFS[16'h1AF4] = 8'h02;
DFS[16'h1AF5] = 8'h85;
DFS[16'h1AF6] = 8'hCA;
DFS[16'h1AF7] = 8'hA9;
DFS[16'h1AF8] = 8'h00;
DFS[16'h1AF9] = 8'h85;
DFS[16'h1AFA] = 8'hCB;
DFS[16'h1AFB] = 8'hA4;
DFS[16'h1AFC] = 8'hCC;
DFS[16'h1AFD] = 8'h20;
DFS[16'h1AFE] = 8'h19;
DFS[16'h1AFF] = 8'h82;
DFS[16'h1B00] = 8'hC0;
DFS[16'h1B01] = 8'hF8;
DFS[16'h1B02] = 8'hD0;
DFS[16'h1B03] = 8'h3C;
DFS[16'h1B04] = 8'h20;
DFS[16'h1B05] = 8'h65;
DFS[16'h1B06] = 8'h80;
DFS[16'h1B07] = 8'h44;
DFS[16'h1B08] = 8'h69;
DFS[16'h1B09] = 8'h73;
DFS[16'h1B0A] = 8'h6B;
DFS[16'h1B0B] = 8'h20;
DFS[16'h1B0C] = 8'h63;
DFS[16'h1B0D] = 8'h6F;
DFS[16'h1B0E] = 8'h6D;
DFS[16'h1B0F] = 8'h70;
DFS[16'h1B10] = 8'h61;
DFS[16'h1B11] = 8'h63;
DFS[16'h1B12] = 8'h74;
DFS[16'h1B13] = 8'h65;
DFS[16'h1B14] = 8'h64;
DFS[16'h1B15] = 8'h20;
DFS[16'h1B16] = 8'hEA;
DFS[16'h1B17] = 8'h38;
DFS[16'h1B18] = 8'hAD;
DFS[16'h1B19] = 8'h07;
DFS[16'h1B1A] = 8'h0F;
DFS[16'h1B1B] = 8'hE5;
DFS[16'h1B1C] = 8'hCA;
DFS[16'h1B1D] = 8'h48;
DFS[16'h1B1E] = 8'hAD;
DFS[16'h1B1F] = 8'h06;
DFS[16'h1B20] = 8'h0F;
DFS[16'h1B21] = 8'h29;
DFS[16'h1B22] = 8'h03;
DFS[16'h1B23] = 8'hE5;
DFS[16'h1B24] = 8'hCB;
DFS[16'h1B25] = 8'h20;
DFS[16'h1B26] = 8'hCA;
DFS[16'h1B27] = 8'h80;
DFS[16'h1B28] = 8'h68;
DFS[16'h1B29] = 8'h20;
DFS[16'h1B2A] = 8'hC2;
DFS[16'h1B2B] = 8'h80;
DFS[16'h1B2C] = 8'h20;
DFS[16'h1B2D] = 8'h65;
DFS[16'h1B2E] = 8'h80;
DFS[16'h1B2F] = 8'h20;
DFS[16'h1B30] = 8'h66;
DFS[16'h1B31] = 8'h72;
DFS[16'h1B32] = 8'h65;
DFS[16'h1B33] = 8'h65;
DFS[16'h1B34] = 8'h20;
DFS[16'h1B35] = 8'h73;
DFS[16'h1B36] = 8'h65;
DFS[16'h1B37] = 8'h63;
DFS[16'h1B38] = 8'h74;
DFS[16'h1B39] = 8'h6F;
DFS[16'h1B3A] = 8'h72;
DFS[16'h1B3B] = 8'h73;
DFS[16'h1B3C] = 8'h0D;
DFS[16'h1B3D] = 8'hA9;
DFS[16'h1B3E] = 8'h04;
DFS[16'h1B3F] = 8'h60;
DFS[16'h1B40] = 8'h84;
DFS[16'h1B41] = 8'hCC;
DFS[16'h1B42] = 8'h20;
DFS[16'h1B43] = 8'hFC;
DFS[16'h1B44] = 8'h82;
DFS[16'h1B45] = 8'hA4;
DFS[16'h1B46] = 8'hCC;
DFS[16'h1B47] = 8'hB9;
DFS[16'h1B48] = 8'h0E;
DFS[16'h1B49] = 8'h0F;
DFS[16'h1B4A] = 8'h29;
DFS[16'h1B4B] = 8'h30;
DFS[16'h1B4C] = 8'h19;
DFS[16'h1B4D] = 8'h0D;
DFS[16'h1B4E] = 8'h0F;
DFS[16'h1B4F] = 8'h19;
DFS[16'h1B50] = 8'h0C;
DFS[16'h1B51] = 8'h0F;
DFS[16'h1B52] = 8'hF0;
DFS[16'h1B53] = 8'h61;
DFS[16'h1B54] = 8'hA9;
DFS[16'h1B55] = 8'h00;
DFS[16'h1B56] = 8'h85;
DFS[16'h1B57] = 8'hBE;
DFS[16'h1B58] = 8'h85;
DFS[16'h1B59] = 8'hC2;
DFS[16'h1B5A] = 8'hA9;
DFS[16'h1B5B] = 8'hFF;
DFS[16'h1B5C] = 8'h18;
DFS[16'h1B5D] = 8'h79;
DFS[16'h1B5E] = 8'h0C;
DFS[16'h1B5F] = 8'h0F;
DFS[16'h1B60] = 8'hA9;
DFS[16'h1B61] = 8'h00;
DFS[16'h1B62] = 8'h79;
DFS[16'h1B63] = 8'h0D;
DFS[16'h1B64] = 8'h0F;
DFS[16'h1B65] = 8'h85;
DFS[16'h1B66] = 8'hC6;
DFS[16'h1B67] = 8'hB9;
DFS[16'h1B68] = 8'h0E;
DFS[16'h1B69] = 8'h0F;
DFS[16'h1B6A] = 8'h08;
DFS[16'h1B6B] = 8'h20;
DFS[16'h1B6C] = 8'hFD;
DFS[16'h1B6D] = 8'h81;
DFS[16'h1B6E] = 8'h28;
DFS[16'h1B6F] = 8'h69;
DFS[16'h1B70] = 8'h00;
DFS[16'h1B71] = 8'h85;
DFS[16'h1B72] = 8'hC7;
DFS[16'h1B73] = 8'hB9;
DFS[16'h1B74] = 8'h0F;
DFS[16'h1B75] = 8'h0F;
DFS[16'h1B76] = 8'h85;
DFS[16'h1B77] = 8'hC8;
DFS[16'h1B78] = 8'hB9;
DFS[16'h1B79] = 8'h0E;
DFS[16'h1B7A] = 8'h0F;
DFS[16'h1B7B] = 8'h29;
DFS[16'h1B7C] = 8'h03;
DFS[16'h1B7D] = 8'h85;
DFS[16'h1B7E] = 8'hC9;
DFS[16'h1B7F] = 8'hC5;
DFS[16'h1B80] = 8'hCB;
DFS[16'h1B81] = 8'hD0;
DFS[16'h1B82] = 8'h14;
DFS[16'h1B83] = 8'hA5;
DFS[16'h1B84] = 8'hC8;
DFS[16'h1B85] = 8'hC5;
DFS[16'h1B86] = 8'hCA;
DFS[16'h1B87] = 8'hD0;
DFS[16'h1B88] = 8'h0E;
DFS[16'h1B89] = 8'h18;
DFS[16'h1B8A] = 8'h65;
DFS[16'h1B8B] = 8'hC6;
DFS[16'h1B8C] = 8'h85;
DFS[16'h1B8D] = 8'hCA;
DFS[16'h1B8E] = 8'hA5;
DFS[16'h1B8F] = 8'hCB;
DFS[16'h1B90] = 8'h65;
DFS[16'h1B91] = 8'hC7;
DFS[16'h1B92] = 8'h85;
DFS[16'h1B93] = 8'hCB;
DFS[16'h1B94] = 8'h4C;
DFS[16'h1B95] = 8'hB5;
DFS[16'h1B96] = 8'h9B;
DFS[16'h1B97] = 8'hA5;
DFS[16'h1B98] = 8'hCA;
DFS[16'h1B99] = 8'h99;
DFS[16'h1B9A] = 8'h0F;
DFS[16'h1B9B] = 8'h0F;
DFS[16'h1B9C] = 8'hB9;
DFS[16'h1B9D] = 8'h0E;
DFS[16'h1B9E] = 8'h0F;
DFS[16'h1B9F] = 8'h29;
DFS[16'h1BA0] = 8'hFC;
DFS[16'h1BA1] = 8'h05;
DFS[16'h1BA2] = 8'hCB;
DFS[16'h1BA3] = 8'h99;
DFS[16'h1BA4] = 8'h0E;
DFS[16'h1BA5] = 8'h0F;
DFS[16'h1BA6] = 8'hA9;
DFS[16'h1BA7] = 8'h00;
DFS[16'h1BA8] = 8'h85;
DFS[16'h1BA9] = 8'hA8;
DFS[16'h1BAA] = 8'h85;
DFS[16'h1BAB] = 8'hA9;
DFS[16'h1BAC] = 8'h20;
DFS[16'h1BAD] = 8'hB4;
DFS[16'h1BAE] = 8'h8A;
DFS[16'h1BAF] = 8'h20;
DFS[16'h1BB0] = 8'h06;
DFS[16'h1BB1] = 8'h9E;
DFS[16'h1BB2] = 8'h20;
DFS[16'h1BB3] = 8'h47;
DFS[16'h1BB4] = 8'h83;
DFS[16'h1BB5] = 8'hA4;
DFS[16'h1BB6] = 8'hCC;
DFS[16'h1BB7] = 8'h20;
DFS[16'h1BB8] = 8'h01;
DFS[16'h1BB9] = 8'h83;
DFS[16'h1BBA] = 8'h4C;
DFS[16'h1BBB] = 8'hFB;
DFS[16'h1BBC] = 8'h9A;
DFS[16'h1BBD] = 8'h2C;
DFS[16'h1BBE] = 8'hC8;
DFS[16'h1BBF] = 8'h10;
DFS[16'h1BC0] = 8'h10;
DFS[16'h1BC1] = 8'h75;
DFS[16'h1BC2] = 8'h20;
DFS[16'h1BC3] = 8'h33;
DFS[16'h1BC4] = 8'h80;
DFS[16'h1BC5] = 8'hBD;
DFS[16'h1BC6] = 8'h4E;
DFS[16'h1BC7] = 8'h6F;
DFS[16'h1BC8] = 8'h74;
DFS[16'h1BC9] = 8'h20;
DFS[16'h1BCA] = 8'h65;
DFS[16'h1BCB] = 8'h6E;
DFS[16'h1BCC] = 8'h61;
DFS[16'h1BCD] = 8'h62;
DFS[16'h1BCE] = 8'h6C;
DFS[16'h1BCF] = 8'h65;
DFS[16'h1BD0] = 8'h64;
DFS[16'h1BD1] = 8'h00;
DFS[16'h1BD2] = 8'h20;
DFS[16'h1BD3] = 8'hBF;
DFS[16'h1BD4] = 8'h86;
DFS[16'h1BD5] = 8'hD0;
DFS[16'h1BD6] = 8'h03;
DFS[16'h1BD7] = 8'h4C;
DFS[16'h1BD8] = 8'h06;
DFS[16'h1BD9] = 8'h9A;
DFS[16'h1BDA] = 8'h20;
DFS[16'h1BDB] = 8'h5D;
DFS[16'h1BDC] = 8'h83;
DFS[16'h1BDD] = 8'h8D;
DFS[16'h1BDE] = 8'hD2;
DFS[16'h1BDF] = 8'h10;
DFS[16'h1BE0] = 8'h20;
DFS[16'h1BE1] = 8'hBF;
DFS[16'h1BE2] = 8'h86;
DFS[16'h1BE3] = 8'hF0;
DFS[16'h1BE4] = 8'hF2;
DFS[16'h1BE5] = 8'h20;
DFS[16'h1BE6] = 8'h5D;
DFS[16'h1BE7] = 8'h83;
DFS[16'h1BE8] = 8'h8D;
DFS[16'h1BE9] = 8'hD3;
DFS[16'h1BEA] = 8'h10;
DFS[16'h1BEB] = 8'h98;
DFS[16'h1BEC] = 8'h48;
DFS[16'h1BED] = 8'hA9;
DFS[16'h1BEE] = 8'h00;
DFS[16'h1BEF] = 8'h85;
DFS[16'h1BF0] = 8'hA9;
DFS[16'h1BF1] = 8'hAD;
DFS[16'h1BF2] = 8'hD3;
DFS[16'h1BF3] = 8'h10;
DFS[16'h1BF4] = 8'hCD;
DFS[16'h1BF5] = 8'hD2;
DFS[16'h1BF6] = 8'h10;
DFS[16'h1BF7] = 8'hD0;
DFS[16'h1BF8] = 8'h06;
DFS[16'h1BF9] = 8'hA9;
DFS[16'h1BFA] = 8'hFF;
DFS[16'h1BFB] = 8'h85;
DFS[16'h1BFC] = 8'hA9;
DFS[16'h1BFD] = 8'h85;
DFS[16'h1BFE] = 8'hAA;
DFS[16'h1BFF] = 8'h20;
DFS[16'h1C00] = 8'h79;
DFS[16'h1C01] = 8'h98;
DFS[16'h1C02] = 8'h20;
DFS[16'h1C03] = 8'h65;
DFS[16'h1C04] = 8'h80;
DFS[16'h1C05] = 8'h43;
DFS[16'h1C06] = 8'h6F;
DFS[16'h1C07] = 8'h70;
DFS[16'h1C08] = 8'h79;
DFS[16'h1C09] = 8'h69;
DFS[16'h1C0A] = 8'h6E;
DFS[16'h1C0B] = 8'h67;
DFS[16'h1C0C] = 8'h20;
DFS[16'h1C0D] = 8'h66;
DFS[16'h1C0E] = 8'h72;
DFS[16'h1C0F] = 8'h6F;
DFS[16'h1C10] = 8'h6D;
DFS[16'h1C11] = 8'h20;
DFS[16'h1C12] = 8'h64;
DFS[16'h1C13] = 8'h72;
DFS[16'h1C14] = 8'h69;
DFS[16'h1C15] = 8'h76;
DFS[16'h1C16] = 8'h65;
DFS[16'h1C17] = 8'h20;
DFS[16'h1C18] = 8'hAD;
DFS[16'h1C19] = 8'hD2;
DFS[16'h1C1A] = 8'h10;
DFS[16'h1C1B] = 8'h20;
DFS[16'h1C1C] = 8'hCA;
DFS[16'h1C1D] = 8'h80;
DFS[16'h1C1E] = 8'h20;
DFS[16'h1C1F] = 8'h65;
DFS[16'h1C20] = 8'h80;
DFS[16'h1C21] = 8'h20;
DFS[16'h1C22] = 8'h74;
DFS[16'h1C23] = 8'h6F;
DFS[16'h1C24] = 8'h20;
DFS[16'h1C25] = 8'h64;
DFS[16'h1C26] = 8'h72;
DFS[16'h1C27] = 8'h69;
DFS[16'h1C28] = 8'h76;
DFS[16'h1C29] = 8'h65;
DFS[16'h1C2A] = 8'h20;
DFS[16'h1C2B] = 8'hAD;
DFS[16'h1C2C] = 8'hD3;
DFS[16'h1C2D] = 8'h10;
DFS[16'h1C2E] = 8'h20;
DFS[16'h1C2F] = 8'hCA;
DFS[16'h1C30] = 8'h80;
DFS[16'h1C31] = 8'h20;
DFS[16'h1C32] = 8'h9A;
DFS[16'h1C33] = 8'h9F;
DFS[16'h1C34] = 8'h68;
DFS[16'h1C35] = 8'hA8;
DFS[16'h1C36] = 8'h18;
DFS[16'h1C37] = 8'h60;
DFS[16'h1C38] = 8'h20;
DFS[16'h1C39] = 8'hE1;
DFS[16'h1C3A] = 8'h83;
DFS[16'h1C3B] = 8'h24;
DFS[16'h1C3C] = 8'hA9;
DFS[16'h1C3D] = 8'h10;
DFS[16'h1C3E] = 8'h0B;
DFS[16'h1C3F] = 8'hA9;
DFS[16'h1C40] = 8'h00;
DFS[16'h1C41] = 8'hF0;
DFS[16'h1C42] = 8'h0A;
DFS[16'h1C43] = 8'h20;
DFS[16'h1C44] = 8'hE1;
DFS[16'h1C45] = 8'h83;
DFS[16'h1C46] = 8'h24;
DFS[16'h1C47] = 8'hA9;
DFS[16'h1C48] = 8'h30;
DFS[16'h1C49] = 8'h01;
DFS[16'h1C4A] = 8'h60;
DFS[16'h1C4B] = 8'hA9;
DFS[16'h1C4C] = 8'h80;
DFS[16'h1C4D] = 8'hC5;
DFS[16'h1C4E] = 8'hAA;
DFS[16'h1C4F] = 8'hF0;
DFS[16'h1C50] = 8'hF9;
DFS[16'h1C51] = 8'h85;
DFS[16'h1C52] = 8'hAA;
DFS[16'h1C53] = 8'h20;
DFS[16'h1C54] = 8'h65;
DFS[16'h1C55] = 8'h80;
DFS[16'h1C56] = 8'h49;
DFS[16'h1C57] = 8'h6E;
DFS[16'h1C58] = 8'h73;
DFS[16'h1C59] = 8'h65;
DFS[16'h1C5A] = 8'h72;
DFS[16'h1C5B] = 8'h74;
DFS[16'h1C5C] = 8'h20;
DFS[16'h1C5D] = 8'hEA;
DFS[16'h1C5E] = 8'h24;
DFS[16'h1C5F] = 8'hAA;
DFS[16'h1C60] = 8'h30;
DFS[16'h1C61] = 8'h0B;
DFS[16'h1C62] = 8'h20;
DFS[16'h1C63] = 8'h65;
DFS[16'h1C64] = 8'h80;
DFS[16'h1C65] = 8'h73;
DFS[16'h1C66] = 8'h6F;
DFS[16'h1C67] = 8'h75;
DFS[16'h1C68] = 8'h72;
DFS[16'h1C69] = 8'h63;
DFS[16'h1C6A] = 8'h65;
DFS[16'h1C6B] = 8'h90;
DFS[16'h1C6C] = 8'h0F;
DFS[16'h1C6D] = 8'h20;
DFS[16'h1C6E] = 8'h65;
DFS[16'h1C6F] = 8'h80;
DFS[16'h1C70] = 8'h64;
DFS[16'h1C71] = 8'h65;
DFS[16'h1C72] = 8'h73;
DFS[16'h1C73] = 8'h74;
DFS[16'h1C74] = 8'h69;
DFS[16'h1C75] = 8'h6E;
DFS[16'h1C76] = 8'h61;
DFS[16'h1C77] = 8'h74;
DFS[16'h1C78] = 8'h69;
DFS[16'h1C79] = 8'h6F;
DFS[16'h1C7A] = 8'h6E;
DFS[16'h1C7B] = 8'hEA;
DFS[16'h1C7C] = 8'h20;
DFS[16'h1C7D] = 8'h65;
DFS[16'h1C7E] = 8'h80;
DFS[16'h1C7F] = 8'h20;
DFS[16'h1C80] = 8'h64;
DFS[16'h1C81] = 8'h69;
DFS[16'h1C82] = 8'h73;
DFS[16'h1C83] = 8'h6B;
DFS[16'h1C84] = 8'h20;
DFS[16'h1C85] = 8'h61;
DFS[16'h1C86] = 8'h6E;
DFS[16'h1C87] = 8'h64;
DFS[16'h1C88] = 8'h20;
DFS[16'h1C89] = 8'h68;
DFS[16'h1C8A] = 8'h69;
DFS[16'h1C8B] = 8'h74;
DFS[16'h1C8C] = 8'h20;
DFS[16'h1C8D] = 8'h61;
DFS[16'h1C8E] = 8'h20;
DFS[16'h1C8F] = 8'h6B;
DFS[16'h1C90] = 8'h65;
DFS[16'h1C91] = 8'h79;
DFS[16'h1C92] = 8'hEA;
DFS[16'h1C93] = 8'h20;
DFS[16'h1C94] = 8'h06;
DFS[16'h1C95] = 8'h99;
DFS[16'h1C96] = 8'h20;
DFS[16'h1C97] = 8'hE0;
DFS[16'h1C98] = 8'hFF;
DFS[16'h1C99] = 8'hB0;
DFS[16'h1C9A] = 8'h19;
DFS[16'h1C9B] = 8'h4C;
DFS[16'h1C9C] = 8'h9A;
DFS[16'h1C9D] = 8'h9F;
DFS[16'h1C9E] = 8'h20;
DFS[16'h1C9F] = 8'h06;
DFS[16'h1CA0] = 8'h99;
DFS[16'h1CA1] = 8'h20;
DFS[16'h1CA2] = 8'hE0;
DFS[16'h1CA3] = 8'hFF;
DFS[16'h1CA4] = 8'hB0;
DFS[16'h1CA5] = 8'h0E;
DFS[16'h1CA6] = 8'h29;
DFS[16'h1CA7] = 8'h5F;
DFS[16'h1CA8] = 8'hC9;
DFS[16'h1CA9] = 8'h59;
DFS[16'h1CAA] = 8'h08;
DFS[16'h1CAB] = 8'hF0;
DFS[16'h1CAC] = 8'h02;
DFS[16'h1CAD] = 8'hA9;
DFS[16'h1CAE] = 8'h4E;
DFS[16'h1CAF] = 8'h20;
DFS[16'h1CB0] = 8'h9C;
DFS[16'h1CB1] = 8'h80;
DFS[16'h1CB2] = 8'h28;
DFS[16'h1CB3] = 8'h60;
DFS[16'h1CB4] = 8'hA6;
DFS[16'h1CB5] = 8'hB6;
DFS[16'h1CB6] = 8'h9A;
DFS[16'h1CB7] = 8'h60;
DFS[16'h1CB8] = 8'h4C;
DFS[16'h1CB9] = 8'h58;
DFS[16'h1CBA] = 8'h89;
DFS[16'h1CBB] = 8'h20;
DFS[16'h1CBC] = 8'hBD;
DFS[16'h1CBD] = 8'h9B;
DFS[16'h1CBE] = 8'h20;
DFS[16'h1CBF] = 8'hD2;
DFS[16'h1CC0] = 8'h9B;
DFS[16'h1CC1] = 8'hA9;
DFS[16'h1CC2] = 8'h00;
DFS[16'h1CC3] = 8'h85;
DFS[16'h1CC4] = 8'hC9;
DFS[16'h1CC5] = 8'h85;
DFS[16'h1CC6] = 8'hCB;
DFS[16'h1CC7] = 8'h85;
DFS[16'h1CC8] = 8'hCA;
DFS[16'h1CC9] = 8'h85;
DFS[16'h1CCA] = 8'hC8;
DFS[16'h1CCB] = 8'h85;
DFS[16'h1CCC] = 8'hA8;
DFS[16'h1CCD] = 8'h20;
DFS[16'h1CCE] = 8'h38;
DFS[16'h1CCF] = 8'h9C;
DFS[16'h1CD0] = 8'hAD;
DFS[16'h1CD1] = 8'hD2;
DFS[16'h1CD2] = 8'h10;
DFS[16'h1CD3] = 8'h85;
DFS[16'h1CD4] = 8'hCF;
DFS[16'h1CD5] = 8'h20;
DFS[16'h1CD6] = 8'h4D;
DFS[16'h1CD7] = 8'hAB;
DFS[16'h1CD8] = 8'hAD;
DFS[16'h1CD9] = 8'h07;
DFS[16'h1CDA] = 8'h0F;
DFS[16'h1CDB] = 8'h85;
DFS[16'h1CDC] = 8'hC6;
DFS[16'h1CDD] = 8'hAD;
DFS[16'h1CDE] = 8'h06;
DFS[16'h1CDF] = 8'h0F;
DFS[16'h1CE0] = 8'h29;
DFS[16'h1CE1] = 8'h03;
DFS[16'h1CE2] = 8'h85;
DFS[16'h1CE3] = 8'hC7;
DFS[16'h1CE4] = 8'hAD;
DFS[16'h1CE5] = 8'h06;
DFS[16'h1CE6] = 8'h0F;
DFS[16'h1CE7] = 8'h29;
DFS[16'h1CE8] = 8'hF0;
DFS[16'h1CE9] = 8'h8D;
DFS[16'h1CEA] = 8'hD8;
DFS[16'h1CEB] = 8'h10;
DFS[16'h1CEC] = 8'h20;
DFS[16'h1CED] = 8'h43;
DFS[16'h1CEE] = 8'h9C;
DFS[16'h1CEF] = 8'hAD;
DFS[16'h1CF0] = 8'hD3;
DFS[16'h1CF1] = 8'h10;
DFS[16'h1CF2] = 8'h85;
DFS[16'h1CF3] = 8'hCF;
DFS[16'h1CF4] = 8'h20;
DFS[16'h1CF5] = 8'h4D;
DFS[16'h1CF6] = 8'hAB;
DFS[16'h1CF7] = 8'hAD;
DFS[16'h1CF8] = 8'h06;
DFS[16'h1CF9] = 8'h0F;
DFS[16'h1CFA] = 8'h29;
DFS[16'h1CFB] = 8'h03;
DFS[16'h1CFC] = 8'hC5;
DFS[16'h1CFD] = 8'hC7;
DFS[16'h1CFE] = 8'h90;
DFS[16'h1CFF] = 8'hB8;
DFS[16'h1D00] = 8'hD0;
DFS[16'h1D01] = 8'h07;
DFS[16'h1D02] = 8'hAD;
DFS[16'h1D03] = 8'h07;
DFS[16'h1D04] = 8'h0F;
DFS[16'h1D05] = 8'hC5;
DFS[16'h1D06] = 8'hC6;
DFS[16'h1D07] = 8'h90;
DFS[16'h1D08] = 8'hAF;
DFS[16'h1D09] = 8'h20;
DFS[16'h1D0A] = 8'h06;
DFS[16'h1D0B] = 8'h9E;
DFS[16'h1D0C] = 8'hAD;
DFS[16'h1D0D] = 8'h06;
DFS[16'h1D0E] = 8'h0F;
DFS[16'h1D0F] = 8'h48;
DFS[16'h1D10] = 8'hAD;
DFS[16'h1D11] = 8'h07;
DFS[16'h1D12] = 8'h0F;
DFS[16'h1D13] = 8'h48;
DFS[16'h1D14] = 8'h20;
DFS[16'h1D15] = 8'h4D;
DFS[16'h1D16] = 8'hAB;
DFS[16'h1D17] = 8'h68;
DFS[16'h1D18] = 8'h8D;
DFS[16'h1D19] = 8'h07;
DFS[16'h1D1A] = 8'h0F;
DFS[16'h1D1B] = 8'h68;
DFS[16'h1D1C] = 8'h29;
DFS[16'h1D1D] = 8'h0F;
DFS[16'h1D1E] = 8'h0D;
DFS[16'h1D1F] = 8'hD8;
DFS[16'h1D20] = 8'h10;
DFS[16'h1D21] = 8'h8D;
DFS[16'h1D22] = 8'h06;
DFS[16'h1D23] = 8'h0F;
DFS[16'h1D24] = 8'h4C;
DFS[16'h1D25] = 8'hB4;
DFS[16'h1D26] = 8'h8A;
DFS[16'h1D27] = 8'h20;
DFS[16'h1D28] = 8'h5E;
DFS[16'h1D29] = 8'h82;
DFS[16'h1D2A] = 8'h20;
DFS[16'h1D2B] = 8'hD2;
DFS[16'h1D2C] = 8'h9B;
DFS[16'h1D2D] = 8'h20;
DFS[16'h1D2E] = 8'hBF;
DFS[16'h1D2F] = 8'h86;
DFS[16'h1D30] = 8'hD0;
DFS[16'h1D31] = 8'h03;
DFS[16'h1D32] = 8'h4C;
DFS[16'h1D33] = 8'h06;
DFS[16'h1D34] = 8'h9A;
DFS[16'h1D35] = 8'h20;
DFS[16'h1D36] = 8'hFE;
DFS[16'h1D37] = 8'h80;
DFS[16'h1D38] = 8'h20;
DFS[16'h1D39] = 8'h38;
DFS[16'h1D3A] = 8'h9C;
DFS[16'h1D3B] = 8'hAD;
DFS[16'h1D3C] = 8'hD2;
DFS[16'h1D3D] = 8'h10;
DFS[16'h1D3E] = 8'h20;
DFS[16'h1D3F] = 8'h7E;
DFS[16'h1D40] = 8'h87;
DFS[16'h1D41] = 8'h20;
DFS[16'h1D42] = 8'h96;
DFS[16'h1D43] = 8'h82;
DFS[16'h1D44] = 8'hB0;
DFS[16'h1D45] = 8'h03;
DFS[16'h1D46] = 8'h4C;
DFS[16'h1D47] = 8'h76;
DFS[16'h1D48] = 8'h82;
DFS[16'h1D49] = 8'h84;
DFS[16'h1D4A] = 8'hAB;
DFS[16'h1D4B] = 8'h20;
DFS[16'h1D4C] = 8'h01;
DFS[16'h1D4D] = 8'h83;
DFS[16'h1D4E] = 8'hA2;
DFS[16'h1D4F] = 8'h00;
DFS[16'h1D50] = 8'hB5;
DFS[16'h1D51] = 8'hC7;
DFS[16'h1D52] = 8'h9D;
DFS[16'h1D53] = 8'h58;
DFS[16'h1D54] = 8'h10;
DFS[16'h1D55] = 8'hB9;
DFS[16'h1D56] = 8'h08;
DFS[16'h1D57] = 8'h0E;
DFS[16'h1D58] = 8'h95;
DFS[16'h1D59] = 8'hC7;
DFS[16'h1D5A] = 8'h9D;
DFS[16'h1D5B] = 8'h50;
DFS[16'h1D5C] = 8'h10;
DFS[16'h1D5D] = 8'hB9;
DFS[16'h1D5E] = 8'h08;
DFS[16'h1D5F] = 8'h0F;
DFS[16'h1D60] = 8'h95;
DFS[16'h1D61] = 8'hBD;
DFS[16'h1D62] = 8'h9D;
DFS[16'h1D63] = 8'h47;
DFS[16'h1D64] = 8'h10;
DFS[16'h1D65] = 8'hE8;
DFS[16'h1D66] = 8'hC8;
DFS[16'h1D67] = 8'hE0;
DFS[16'h1D68] = 8'h08;
DFS[16'h1D69] = 8'hD0;
DFS[16'h1D6A] = 8'hE5;
DFS[16'h1D6B] = 8'hA5;
DFS[16'h1D6C] = 8'hC3;
DFS[16'h1D6D] = 8'h20;
DFS[16'h1D6E] = 8'hFD;
DFS[16'h1D6F] = 8'h81;
DFS[16'h1D70] = 8'h85;
DFS[16'h1D71] = 8'hC5;
DFS[16'h1D72] = 8'hA5;
DFS[16'h1D73] = 8'hC1;
DFS[16'h1D74] = 8'h18;
DFS[16'h1D75] = 8'h69;
DFS[16'h1D76] = 8'hFF;
DFS[16'h1D77] = 8'hA5;
DFS[16'h1D78] = 8'hC2;
DFS[16'h1D79] = 8'h69;
DFS[16'h1D7A] = 8'h00;
DFS[16'h1D7B] = 8'h85;
DFS[16'h1D7C] = 8'hC6;
DFS[16'h1D7D] = 8'hA5;
DFS[16'h1D7E] = 8'hC5;
DFS[16'h1D7F] = 8'h69;
DFS[16'h1D80] = 8'h00;
DFS[16'h1D81] = 8'h85;
DFS[16'h1D82] = 8'hC7;
DFS[16'h1D83] = 8'hAD;
DFS[16'h1D84] = 8'h4E;
DFS[16'h1D85] = 8'h10;
DFS[16'h1D86] = 8'h85;
DFS[16'h1D87] = 8'hC8;
DFS[16'h1D88] = 8'hAD;
DFS[16'h1D89] = 8'h4D;
DFS[16'h1D8A] = 8'h10;
DFS[16'h1D8B] = 8'h29;
DFS[16'h1D8C] = 8'h03;
DFS[16'h1D8D] = 8'h85;
DFS[16'h1D8E] = 8'hC9;
DFS[16'h1D8F] = 8'hA9;
DFS[16'h1D90] = 8'hFF;
DFS[16'h1D91] = 8'h85;
DFS[16'h1D92] = 8'hA8;
DFS[16'h1D93] = 8'h20;
DFS[16'h1D94] = 8'h06;
DFS[16'h1D95] = 8'h9E;
DFS[16'h1D96] = 8'h20;
DFS[16'h1D97] = 8'h38;
DFS[16'h1D98] = 8'h9C;
DFS[16'h1D99] = 8'hAD;
DFS[16'h1D9A] = 8'hD2;
DFS[16'h1D9B] = 8'h10;
DFS[16'h1D9C] = 8'h20;
DFS[16'h1D9D] = 8'h7E;
DFS[16'h1D9E] = 8'h87;
DFS[16'h1D9F] = 8'h20;
DFS[16'h1DA0] = 8'h47;
DFS[16'h1DA1] = 8'h83;
DFS[16'h1DA2] = 8'hA2;
DFS[16'h1DA3] = 8'h07;
DFS[16'h1DA4] = 8'hBD;
DFS[16'h1DA5] = 8'h58;
DFS[16'h1DA6] = 8'h10;
DFS[16'h1DA7] = 8'h95;
DFS[16'h1DA8] = 8'hC7;
DFS[16'h1DA9] = 8'hCA;
DFS[16'h1DAA] = 8'h10;
DFS[16'h1DAB] = 8'hF8;
DFS[16'h1DAC] = 8'hA4;
DFS[16'h1DAD] = 8'hAB;
DFS[16'h1DAE] = 8'h8C;
DFS[16'h1DAF] = 8'hCE;
DFS[16'h1DB0] = 8'h10;
DFS[16'h1DB1] = 8'h20;
DFS[16'h1DB2] = 8'h9D;
DFS[16'h1DB3] = 8'h82;
DFS[16'h1DB4] = 8'hB0;
DFS[16'h1DB5] = 8'h93;
DFS[16'h1DB6] = 8'h60;
DFS[16'h1DB7] = 8'h20;
DFS[16'h1DB8] = 8'hF5;
DFS[16'h1DB9] = 8'h9D;
DFS[16'h1DBA] = 8'h20;
DFS[16'h1DBB] = 8'h43;
DFS[16'h1DBC] = 8'h9C;
DFS[16'h1DBD] = 8'hAD;
DFS[16'h1DBE] = 8'hD3;
DFS[16'h1DBF] = 8'h10;
DFS[16'h1DC0] = 8'h85;
DFS[16'h1DC1] = 8'hCF;
DFS[16'h1DC2] = 8'hA5;
DFS[16'h1DC3] = 8'hCE;
DFS[16'h1DC4] = 8'h48;
DFS[16'h1DC5] = 8'h20;
DFS[16'h1DC6] = 8'h47;
DFS[16'h1DC7] = 8'h83;
DFS[16'h1DC8] = 8'h20;
DFS[16'h1DC9] = 8'h96;
DFS[16'h1DCA] = 8'h82;
DFS[16'h1DCB] = 8'h90;
DFS[16'h1DCC] = 8'h03;
DFS[16'h1DCD] = 8'h20;
DFS[16'h1DCE] = 8'hD1;
DFS[16'h1DCF] = 8'h82;
DFS[16'h1DD0] = 8'h68;
DFS[16'h1DD1] = 8'h85;
DFS[16'h1DD2] = 8'hCE;
DFS[16'h1DD3] = 8'h20;
DFS[16'h1DD4] = 8'h3F;
DFS[16'h1DD5] = 8'h8A;
DFS[16'h1DD6] = 8'h20;
DFS[16'h1DD7] = 8'h56;
DFS[16'h1DD8] = 8'h8A;
DFS[16'h1DD9] = 8'hA5;
DFS[16'h1DDA] = 8'hC4;
DFS[16'h1DDB] = 8'h20;
DFS[16'h1DDC] = 8'hFD;
DFS[16'h1DDD] = 8'h81;
DFS[16'h1DDE] = 8'h85;
DFS[16'h1DDF] = 8'hC6;
DFS[16'h1DE0] = 8'h20;
DFS[16'h1DE1] = 8'h9D;
DFS[16'h1DE2] = 8'h89;
DFS[16'h1DE3] = 8'hA5;
DFS[16'h1DE4] = 8'hC4;
DFS[16'h1DE5] = 8'h29;
DFS[16'h1DE6] = 8'h03;
DFS[16'h1DE7] = 8'h48;
DFS[16'h1DE8] = 8'hA5;
DFS[16'h1DE9] = 8'hC5;
DFS[16'h1DEA] = 8'h48;
DFS[16'h1DEB] = 8'h20;
DFS[16'h1DEC] = 8'hF5;
DFS[16'h1DED] = 8'h9D;
DFS[16'h1DEE] = 8'h68;
DFS[16'h1DEF] = 8'h85;
DFS[16'h1DF0] = 8'hCA;
DFS[16'h1DF1] = 8'h68;
DFS[16'h1DF2] = 8'h85;
DFS[16'h1DF3] = 8'hCB;
DFS[16'h1DF4] = 8'h60;
DFS[16'h1DF5] = 8'hA2;
DFS[16'h1DF6] = 8'h11;
DFS[16'h1DF7] = 8'hBD;
DFS[16'h1DF8] = 8'h45;
DFS[16'h1DF9] = 8'h10;
DFS[16'h1DFA] = 8'hB4;
DFS[16'h1DFB] = 8'hBC;
DFS[16'h1DFC] = 8'h95;
DFS[16'h1DFD] = 8'hBC;
DFS[16'h1DFE] = 8'h98;
DFS[16'h1DFF] = 8'h9D;
DFS[16'h1E00] = 8'h45;
DFS[16'h1E01] = 8'h10;
DFS[16'h1E02] = 8'hCA;
DFS[16'h1E03] = 8'h10;
DFS[16'h1E04] = 8'hF2;
DFS[16'h1E05] = 8'h60;
DFS[16'h1E06] = 8'h20;
DFS[16'h1E07] = 8'h8D;
DFS[16'h1E08] = 8'hA0;
DFS[16'h1E09] = 8'hA9;
DFS[16'h1E0A] = 8'h00;
DFS[16'h1E0B] = 8'h85;
DFS[16'h1E0C] = 8'hBE;
DFS[16'h1E0D] = 8'h85;
DFS[16'h1E0E] = 8'hC2;
DFS[16'h1E0F] = 8'hA5;
DFS[16'h1E10] = 8'hC6;
DFS[16'h1E11] = 8'hA8;
DFS[16'h1E12] = 8'hCD;
DFS[16'h1E13] = 8'hD1;
DFS[16'h1E14] = 8'h10;
DFS[16'h1E15] = 8'hA5;
DFS[16'h1E16] = 8'hC7;
DFS[16'h1E17] = 8'hE9;
DFS[16'h1E18] = 8'h00;
DFS[16'h1E19] = 8'h90;
DFS[16'h1E1A] = 8'h03;
DFS[16'h1E1B] = 8'hAC;
DFS[16'h1E1C] = 8'hD1;
DFS[16'h1E1D] = 8'h10;
DFS[16'h1E1E] = 8'h84;
DFS[16'h1E1F] = 8'hC3;
DFS[16'h1E20] = 8'hA5;
DFS[16'h1E21] = 8'hC8;
DFS[16'h1E22] = 8'h85;
DFS[16'h1E23] = 8'hC5;
DFS[16'h1E24] = 8'hA5;
DFS[16'h1E25] = 8'hC9;
DFS[16'h1E26] = 8'h85;
DFS[16'h1E27] = 8'hC4;
DFS[16'h1E28] = 8'hAD;
DFS[16'h1E29] = 8'hD0;
DFS[16'h1E2A] = 8'h10;
DFS[16'h1E2B] = 8'h85;
DFS[16'h1E2C] = 8'hBF;
DFS[16'h1E2D] = 8'hAD;
DFS[16'h1E2E] = 8'hD2;
DFS[16'h1E2F] = 8'h10;
DFS[16'h1E30] = 8'h85;
DFS[16'h1E31] = 8'hCF;
DFS[16'h1E32] = 8'h20;
DFS[16'h1E33] = 8'h38;
DFS[16'h1E34] = 8'h9C;
DFS[16'h1E35] = 8'h20;
DFS[16'h1E36] = 8'h0B;
DFS[16'h1E37] = 8'hB9;
DFS[16'h1E38] = 8'h20;
DFS[16'h1E39] = 8'hC6;
DFS[16'h1E3A] = 8'h87;
DFS[16'h1E3B] = 8'hAD;
DFS[16'h1E3C] = 8'hD3;
DFS[16'h1E3D] = 8'h10;
DFS[16'h1E3E] = 8'h85;
DFS[16'h1E3F] = 8'hCF;
DFS[16'h1E40] = 8'h24;
DFS[16'h1E41] = 8'hA8;
DFS[16'h1E42] = 8'h10;
DFS[16'h1E43] = 8'h07;
DFS[16'h1E44] = 8'h20;
DFS[16'h1E45] = 8'hB7;
DFS[16'h1E46] = 8'h9D;
DFS[16'h1E47] = 8'hA9;
DFS[16'h1E48] = 8'h00;
DFS[16'h1E49] = 8'h85;
DFS[16'h1E4A] = 8'hA8;
DFS[16'h1E4B] = 8'hA5;
DFS[16'h1E4C] = 8'hCA;
DFS[16'h1E4D] = 8'h85;
DFS[16'h1E4E] = 8'hC5;
DFS[16'h1E4F] = 8'hA5;
DFS[16'h1E50] = 8'hCB;
DFS[16'h1E51] = 8'h85;
DFS[16'h1E52] = 8'hC4;
DFS[16'h1E53] = 8'hAD;
DFS[16'h1E54] = 8'hD0;
DFS[16'h1E55] = 8'h10;
DFS[16'h1E56] = 8'h85;
DFS[16'h1E57] = 8'hBF;
DFS[16'h1E58] = 8'h20;
DFS[16'h1E59] = 8'h43;
DFS[16'h1E5A] = 8'h9C;
DFS[16'h1E5B] = 8'h20;
DFS[16'h1E5C] = 8'h0B;
DFS[16'h1E5D] = 8'hB9;
DFS[16'h1E5E] = 8'h20;
DFS[16'h1E5F] = 8'h8F;
DFS[16'h1E60] = 8'h87;
DFS[16'h1E61] = 8'hA5;
DFS[16'h1E62] = 8'hC3;
DFS[16'h1E63] = 8'h18;
DFS[16'h1E64] = 8'h65;
DFS[16'h1E65] = 8'hCA;
DFS[16'h1E66] = 8'h85;
DFS[16'h1E67] = 8'hCA;
DFS[16'h1E68] = 8'h90;
DFS[16'h1E69] = 8'h02;
DFS[16'h1E6A] = 8'hE6;
DFS[16'h1E6B] = 8'hCB;
DFS[16'h1E6C] = 8'hA5;
DFS[16'h1E6D] = 8'hC3;
DFS[16'h1E6E] = 8'h18;
DFS[16'h1E6F] = 8'h65;
DFS[16'h1E70] = 8'hC8;
DFS[16'h1E71] = 8'h85;
DFS[16'h1E72] = 8'hC8;
DFS[16'h1E73] = 8'h90;
DFS[16'h1E74] = 8'h02;
DFS[16'h1E75] = 8'hE6;
DFS[16'h1E76] = 8'hC9;
DFS[16'h1E77] = 8'h38;
DFS[16'h1E78] = 8'hA5;
DFS[16'h1E79] = 8'hC6;
DFS[16'h1E7A] = 8'hE5;
DFS[16'h1E7B] = 8'hC3;
DFS[16'h1E7C] = 8'h85;
DFS[16'h1E7D] = 8'hC6;
DFS[16'h1E7E] = 8'hB0;
DFS[16'h1E7F] = 8'h02;
DFS[16'h1E80] = 8'hC6;
DFS[16'h1E81] = 8'hC7;
DFS[16'h1E82] = 8'h05;
DFS[16'h1E83] = 8'hC7;
DFS[16'h1E84] = 8'hD0;
DFS[16'h1E85] = 8'h89;
DFS[16'h1E86] = 8'h60;
DFS[16'h1E87] = 8'h20;
DFS[16'h1E88] = 8'hD7;
DFS[16'h1E89] = 8'h9F;
DFS[16'h1E8A] = 8'hA9;
DFS[16'h1E8B] = 8'h00;
DFS[16'h1E8C] = 8'hF0;
DFS[16'h1E8D] = 8'h05;
DFS[16'h1E8E] = 8'h20;
DFS[16'h1E8F] = 8'hD7;
DFS[16'h1E90] = 8'h9F;
DFS[16'h1E91] = 8'hA9;
DFS[16'h1E92] = 8'hFF;
DFS[16'h1E93] = 8'h85;
DFS[16'h1E94] = 8'hAB;
DFS[16'h1E95] = 8'hA9;
DFS[16'h1E96] = 8'hC0;
DFS[16'h1E97] = 8'h20;
DFS[16'h1E98] = 8'hCE;
DFS[16'h1E99] = 8'hFF;
DFS[16'h1E9A] = 8'hA8;
DFS[16'h1E9B] = 8'hA9;
DFS[16'h1E9C] = 8'h0D;
DFS[16'h1E9D] = 8'hC0;
DFS[16'h1E9E] = 8'h00;
DFS[16'h1E9F] = 8'hD0;
DFS[16'h1EA0] = 8'h1E;
DFS[16'h1EA1] = 8'h4C;
DFS[16'h1EA2] = 8'h76;
DFS[16'h1EA3] = 8'h82;
DFS[16'h1EA4] = 8'h20;
DFS[16'h1EA5] = 8'hD7;
DFS[16'h1EA6] = 8'hFF;
DFS[16'h1EA7] = 8'hB0;
DFS[16'h1EA8] = 8'h1E;
DFS[16'h1EA9] = 8'hC9;
DFS[16'h1EAA] = 8'h0A;
DFS[16'h1EAB] = 8'hF0;
DFS[16'h1EAC] = 8'hF7;
DFS[16'h1EAD] = 8'h28;
DFS[16'h1EAE] = 8'hD0;
DFS[16'h1EAF] = 8'h08;
DFS[16'h1EB0] = 8'h48;
DFS[16'h1EB1] = 8'h20;
DFS[16'h1EB2] = 8'hA2;
DFS[16'h1EB3] = 8'h9F;
DFS[16'h1EB4] = 8'h20;
DFS[16'h1EB5] = 8'hCE;
DFS[16'h1EB6] = 8'h9F;
DFS[16'h1EB7] = 8'h68;
DFS[16'h1EB8] = 8'h20;
DFS[16'h1EB9] = 8'hE3;
DFS[16'h1EBA] = 8'hFF;
DFS[16'h1EBB] = 8'h24;
DFS[16'h1EBC] = 8'hFF;
DFS[16'h1EBD] = 8'h30;
DFS[16'h1EBE] = 8'h09;
DFS[16'h1EBF] = 8'h25;
DFS[16'h1EC0] = 8'hAB;
DFS[16'h1EC1] = 8'hC9;
DFS[16'h1EC2] = 8'h0D;
DFS[16'h1EC3] = 8'h08;
DFS[16'h1EC4] = 8'h4C;
DFS[16'h1EC5] = 8'hA4;
DFS[16'h1EC6] = 8'h9E;
DFS[16'h1EC7] = 8'h28;
DFS[16'h1EC8] = 8'h20;
DFS[16'h1EC9] = 8'h9A;
DFS[16'h1ECA] = 8'h9F;
DFS[16'h1ECB] = 8'hA9;
DFS[16'h1ECC] = 8'h00;
DFS[16'h1ECD] = 8'h4C;
DFS[16'h1ECE] = 8'hCE;
DFS[16'h1ECF] = 8'hFF;
DFS[16'h1ED0] = 8'h20;
DFS[16'h1ED1] = 8'hD7;
DFS[16'h1ED2] = 8'h9F;
DFS[16'h1ED3] = 8'hA9;
DFS[16'h1ED4] = 8'hC0;
DFS[16'h1ED5] = 8'h20;
DFS[16'h1ED6] = 8'hCE;
DFS[16'h1ED7] = 8'hFF;
DFS[16'h1ED8] = 8'hA8;
DFS[16'h1ED9] = 8'hF0;
DFS[16'h1EDA] = 8'hC6;
DFS[16'h1EDB] = 8'hA6;
DFS[16'h1EDC] = 8'hF4;
DFS[16'h1EDD] = 8'hBD;
DFS[16'h1EDE] = 8'hF0;
DFS[16'h1EDF] = 8'h0D;
DFS[16'h1EE0] = 8'h85;
DFS[16'h1EE1] = 8'hAD;
DFS[16'h1EE2] = 8'hE6;
DFS[16'h1EE3] = 8'hAD;
DFS[16'h1EE4] = 8'h24;
DFS[16'h1EE5] = 8'hFF;
DFS[16'h1EE6] = 8'h30;
DFS[16'h1EE7] = 8'hE3;
DFS[16'h1EE8] = 8'hA5;
DFS[16'h1EE9] = 8'hA9;
DFS[16'h1EEA] = 8'h20;
DFS[16'h1EEB] = 8'hC2;
DFS[16'h1EEC] = 8'h80;
DFS[16'h1EED] = 8'hA5;
DFS[16'h1EEE] = 8'hA8;
DFS[16'h1EEF] = 8'h20;
DFS[16'h1EF0] = 8'hC2;
DFS[16'h1EF1] = 8'h80;
DFS[16'h1EF2] = 8'h20;
DFS[16'h1EF3] = 8'hCE;
DFS[16'h1EF4] = 8'h9F;
DFS[16'h1EF5] = 8'hA9;
DFS[16'h1EF6] = 8'h07;
DFS[16'h1EF7] = 8'h85;
DFS[16'h1EF8] = 8'hAC;
DFS[16'h1EF9] = 8'hA2;
DFS[16'h1EFA] = 8'h00;
DFS[16'h1EFB] = 8'h20;
DFS[16'h1EFC] = 8'hD7;
DFS[16'h1EFD] = 8'hFF;
DFS[16'h1EFE] = 8'hB0;
DFS[16'h1EFF] = 8'h0D;
DFS[16'h1F00] = 8'h81;
DFS[16'h1F01] = 8'hAC;
DFS[16'h1F02] = 8'h20;
DFS[16'h1F03] = 8'hC2;
DFS[16'h1F04] = 8'h80;
DFS[16'h1F05] = 8'h20;
DFS[16'h1F06] = 8'hCE;
DFS[16'h1F07] = 8'h9F;
DFS[16'h1F08] = 8'hC6;
DFS[16'h1F09] = 8'hAC;
DFS[16'h1F0A] = 8'h10;
DFS[16'h1F0B] = 8'hEF;
DFS[16'h1F0C] = 8'h18;
DFS[16'h1F0D] = 8'h08;
DFS[16'h1F0E] = 8'h90;
DFS[16'h1F0F] = 8'h0E;
DFS[16'h1F10] = 8'h20;
DFS[16'h1F11] = 8'h65;
DFS[16'h1F12] = 8'h80;
DFS[16'h1F13] = 8'h2A;
DFS[16'h1F14] = 8'h2A;
DFS[16'h1F15] = 8'h20;
DFS[16'h1F16] = 8'hA9;
DFS[16'h1F17] = 8'h00;
DFS[16'h1F18] = 8'h81;
DFS[16'h1F19] = 8'hAC;
DFS[16'h1F1A] = 8'hC6;
DFS[16'h1F1B] = 8'hAC;
DFS[16'h1F1C] = 8'h10;
DFS[16'h1F1D] = 8'hF2;
DFS[16'h1F1E] = 8'hA9;
DFS[16'h1F1F] = 8'h07;
DFS[16'h1F20] = 8'h85;
DFS[16'h1F21] = 8'hAC;
DFS[16'h1F22] = 8'hA1;
DFS[16'h1F23] = 8'hAC;
DFS[16'h1F24] = 8'hC9;
DFS[16'h1F25] = 8'h7F;
DFS[16'h1F26] = 8'hB0;
DFS[16'h1F27] = 8'h04;
DFS[16'h1F28] = 8'hC9;
DFS[16'h1F29] = 8'h20;
DFS[16'h1F2A] = 8'hB0;
DFS[16'h1F2B] = 8'h02;
DFS[16'h1F2C] = 8'hA9;
DFS[16'h1F2D] = 8'h2E;
DFS[16'h1F2E] = 8'h20;
DFS[16'h1F2F] = 8'hE3;
DFS[16'h1F30] = 8'hFF;
DFS[16'h1F31] = 8'hC6;
DFS[16'h1F32] = 8'hAC;
DFS[16'h1F33] = 8'h10;
DFS[16'h1F34] = 8'hED;
DFS[16'h1F35] = 8'h20;
DFS[16'h1F36] = 8'h9A;
DFS[16'h1F37] = 8'h9F;
DFS[16'h1F38] = 8'hA9;
DFS[16'h1F39] = 8'h08;
DFS[16'h1F3A] = 8'h18;
DFS[16'h1F3B] = 8'h65;
DFS[16'h1F3C] = 8'hA8;
DFS[16'h1F3D] = 8'h85;
DFS[16'h1F3E] = 8'hA8;
DFS[16'h1F3F] = 8'h90;
DFS[16'h1F40] = 8'h02;
DFS[16'h1F41] = 8'hE6;
DFS[16'h1F42] = 8'hA9;
DFS[16'h1F43] = 8'h28;
DFS[16'h1F44] = 8'h90;
DFS[16'h1F45] = 8'h9E;
DFS[16'h1F46] = 8'hB0;
DFS[16'h1F47] = 8'h83;
DFS[16'h1F48] = 8'h20;
DFS[16'h1F49] = 8'hD7;
DFS[16'h1F4A] = 8'h9F;
DFS[16'h1F4B] = 8'hA9;
DFS[16'h1F4C] = 8'h80;
DFS[16'h1F4D] = 8'h20;
DFS[16'h1F4E] = 8'hCE;
DFS[16'h1F4F] = 8'hFF;
DFS[16'h1F50] = 8'h85;
DFS[16'h1F51] = 8'hAB;
DFS[16'h1F52] = 8'h20;
DFS[16'h1F53] = 8'hA2;
DFS[16'h1F54] = 8'h9F;
DFS[16'h1F55] = 8'h20;
DFS[16'h1F56] = 8'hCE;
DFS[16'h1F57] = 8'h9F;
DFS[16'h1F58] = 8'hA6;
DFS[16'h1F59] = 8'hF4;
DFS[16'h1F5A] = 8'hBC;
DFS[16'h1F5B] = 8'hF0;
DFS[16'h1F5C] = 8'h0D;
DFS[16'h1F5D] = 8'hC8;
DFS[16'h1F5E] = 8'h84;
DFS[16'h1F5F] = 8'hAD;
DFS[16'h1F60] = 8'hA2;
DFS[16'h1F61] = 8'hAC;
DFS[16'h1F62] = 8'hA0;
DFS[16'h1F63] = 8'hFF;
DFS[16'h1F64] = 8'h84;
DFS[16'h1F65] = 8'hAE;
DFS[16'h1F66] = 8'h84;
DFS[16'h1F67] = 8'hB0;
DFS[16'h1F68] = 8'hC8;
DFS[16'h1F69] = 8'h84;
DFS[16'h1F6A] = 8'hAC;
DFS[16'h1F6B] = 8'h84;
DFS[16'h1F6C] = 8'hAF;
DFS[16'h1F6D] = 8'h98;
DFS[16'h1F6E] = 8'h20;
DFS[16'h1F6F] = 8'hF1;
DFS[16'h1F70] = 8'hFF;
DFS[16'h1F71] = 8'h08;
DFS[16'h1F72] = 8'h84;
DFS[16'h1F73] = 8'hAA;
DFS[16'h1F74] = 8'hA4;
DFS[16'h1F75] = 8'hAB;
DFS[16'h1F76] = 8'hA2;
DFS[16'h1F77] = 8'h00;
DFS[16'h1F78] = 8'hF0;
DFS[16'h1F79] = 8'h07;
DFS[16'h1F7A] = 8'hA1;
DFS[16'h1F7B] = 8'hAC;
DFS[16'h1F7C] = 8'h20;
DFS[16'h1F7D] = 8'hD4;
DFS[16'h1F7E] = 8'hFF;
DFS[16'h1F7F] = 8'hE6;
DFS[16'h1F80] = 8'hAC;
DFS[16'h1F81] = 8'hA5;
DFS[16'h1F82] = 8'hAC;
DFS[16'h1F83] = 8'hC5;
DFS[16'h1F84] = 8'hAA;
DFS[16'h1F85] = 8'hD0;
DFS[16'h1F86] = 8'hF3;
DFS[16'h1F87] = 8'h28;
DFS[16'h1F88] = 8'hB0;
DFS[16'h1F89] = 8'h08;
DFS[16'h1F8A] = 8'hA9;
DFS[16'h1F8B] = 8'h0D;
DFS[16'h1F8C] = 8'h20;
DFS[16'h1F8D] = 8'hD4;
DFS[16'h1F8E] = 8'hFF;
DFS[16'h1F8F] = 8'h4C;
DFS[16'h1F90] = 8'h52;
DFS[16'h1F91] = 8'h9F;
DFS[16'h1F92] = 8'hA9;
DFS[16'h1F93] = 8'h7E;
DFS[16'h1F94] = 8'h20;
DFS[16'h1F95] = 8'hF4;
DFS[16'h1F96] = 8'hFF;
DFS[16'h1F97] = 8'h20;
DFS[16'h1F98] = 8'hCB;
DFS[16'h1F99] = 8'h9E;
DFS[16'h1F9A] = 8'h48;
DFS[16'h1F9B] = 8'hA9;
DFS[16'h1F9C] = 8'h0D;
DFS[16'h1F9D] = 8'h20;
DFS[16'h1F9E] = 8'h9C;
DFS[16'h1F9F] = 8'h80;
DFS[16'h1FA0] = 8'h68;
DFS[16'h1FA1] = 8'h60;
DFS[16'h1FA2] = 8'hF8;
DFS[16'h1FA3] = 8'h18;
DFS[16'h1FA4] = 8'hA5;
DFS[16'h1FA5] = 8'hA8;
DFS[16'h1FA6] = 8'h69;
DFS[16'h1FA7] = 8'h01;
DFS[16'h1FA8] = 8'h85;
DFS[16'h1FA9] = 8'hA8;
DFS[16'h1FAA] = 8'hA5;
DFS[16'h1FAB] = 8'hA9;
DFS[16'h1FAC] = 8'h69;
DFS[16'h1FAD] = 8'h00;
DFS[16'h1FAE] = 8'h85;
DFS[16'h1FAF] = 8'hA9;
DFS[16'h1FB0] = 8'hD8;
DFS[16'h1FB1] = 8'h18;
DFS[16'h1FB2] = 8'h20;
DFS[16'h1FB3] = 8'hB7;
DFS[16'h1FB4] = 8'h9F;
DFS[16'h1FB5] = 8'hA5;
DFS[16'h1FB6] = 8'hA8;
DFS[16'h1FB7] = 8'h48;
DFS[16'h1FB8] = 8'h08;
DFS[16'h1FB9] = 8'h20;
DFS[16'h1FBA] = 8'h05;
DFS[16'h1FBB] = 8'h82;
DFS[16'h1FBC] = 8'h28;
DFS[16'h1FBD] = 8'h20;
DFS[16'h1FBE] = 8'hC1;
DFS[16'h1FBF] = 8'h9F;
DFS[16'h1FC0] = 8'h68;
DFS[16'h1FC1] = 8'hAA;
DFS[16'h1FC2] = 8'hB0;
DFS[16'h1FC3] = 8'h02;
DFS[16'h1FC4] = 8'hF0;
DFS[16'h1FC5] = 8'h08;
DFS[16'h1FC6] = 8'h20;
DFS[16'h1FC7] = 8'hCA;
DFS[16'h1FC8] = 8'h80;
DFS[16'h1FC9] = 8'h38;
DFS[16'h1FCA] = 8'h60;
DFS[16'h1FCB] = 8'h20;
DFS[16'h1FCC] = 8'hCE;
DFS[16'h1FCD] = 8'h9F;
DFS[16'h1FCE] = 8'h48;
DFS[16'h1FCF] = 8'hA9;
DFS[16'h1FD0] = 8'h20;
DFS[16'h1FD1] = 8'h20;
DFS[16'h1FD2] = 8'h9C;
DFS[16'h1FD3] = 8'h80;
DFS[16'h1FD4] = 8'h68;
DFS[16'h1FD5] = 8'h18;
DFS[16'h1FD6] = 8'h60;
DFS[16'h1FD7] = 8'hBA;
DFS[16'h1FD8] = 8'hA9;
DFS[16'h1FD9] = 8'h00;
DFS[16'h1FDA] = 8'h9D;
DFS[16'h1FDB] = 8'h07;
DFS[16'h1FDC] = 8'h01;
DFS[16'h1FDD] = 8'h88;
DFS[16'h1FDE] = 8'hC8;
DFS[16'h1FDF] = 8'hB1;
DFS[16'h1FE0] = 8'hF2;
DFS[16'h1FE1] = 8'hC9;
DFS[16'h1FE2] = 8'h20;
DFS[16'h1FE3] = 8'hF0;
DFS[16'h1FE4] = 8'hF9;
DFS[16'h1FE5] = 8'hC9;
DFS[16'h1FE6] = 8'h0D;
DFS[16'h1FE7] = 8'hD0;
DFS[16'h1FE8] = 8'h03;
DFS[16'h1FE9] = 8'h4C;
DFS[16'h1FEA] = 8'h06;
DFS[16'h1FEB] = 8'h9A;
DFS[16'h1FEC] = 8'hA9;
DFS[16'h1FED] = 8'h00;
DFS[16'h1FEE] = 8'h85;
DFS[16'h1FEF] = 8'hA8;
DFS[16'h1FF0] = 8'h85;
DFS[16'h1FF1] = 8'hA9;
DFS[16'h1FF2] = 8'h48;
DFS[16'h1FF3] = 8'h98;
DFS[16'h1FF4] = 8'h18;
DFS[16'h1FF5] = 8'h65;
DFS[16'h1FF6] = 8'hF2;
DFS[16'h1FF7] = 8'hAA;
DFS[16'h1FF8] = 8'hA5;
DFS[16'h1FF9] = 8'hF3;
DFS[16'h1FFA] = 8'h69;
DFS[16'h1FFB] = 8'h00;
DFS[16'h1FFC] = 8'hA8;
DFS[16'h1FFD] = 8'h68;
DFS[16'h1FFE] = 8'h60;
DFS[16'h1FFF] = 8'h6D;
DFS[16'h2000] = 8'h20;
DFS[16'h2001] = 8'h7B;
DFS[16'h2002] = 8'hA1;
DFS[16'h2003] = 8'h68;
DFS[16'h2004] = 8'h85;
DFS[16'h2005] = 8'hB8;
DFS[16'h2006] = 8'h68;
DFS[16'h2007] = 8'h85;
DFS[16'h2008] = 8'hB9;
DFS[16'h2009] = 8'h20;
DFS[16'h200A] = 8'h0F;
DFS[16'h200B] = 8'hA0;
DFS[16'h200C] = 8'h4C;
DFS[16'h200D] = 8'h00;
DFS[16'h200E] = 8'h01;
DFS[16'h200F] = 8'hA0;
DFS[16'h2010] = 8'h00;
DFS[16'h2011] = 8'h8C;
DFS[16'h2012] = 8'h00;
DFS[16'h2013] = 8'h01;
DFS[16'h2014] = 8'hC8;
DFS[16'h2015] = 8'hF0;
DFS[16'h2016] = 8'h07;
DFS[16'h2017] = 8'hB1;
DFS[16'h2018] = 8'hB8;
DFS[16'h2019] = 8'h99;
DFS[16'h201A] = 8'h00;
DFS[16'h201B] = 8'h01;
DFS[16'h201C] = 8'hD0;
DFS[16'h201D] = 8'hF6;
DFS[16'h201E] = 8'h60;
DFS[16'h201F] = 8'hA2;
DFS[16'h2020] = 8'hFF;
DFS[16'h2021] = 8'hD0;
DFS[16'h2022] = 8'h02;
DFS[16'h2023] = 8'hA2;
DFS[16'h2024] = 8'h00;
DFS[16'h2025] = 8'hA0;
DFS[16'h2026] = 8'hFF;
DFS[16'h2027] = 8'h8C;
DFS[16'h2028] = 8'h82;
DFS[16'h2029] = 8'h10;
DFS[16'h202A] = 8'h85;
DFS[16'h202B] = 8'hB0;
DFS[16'h202C] = 8'h86;
DFS[16'h202D] = 8'hB1;
DFS[16'h202E] = 8'h8D;
DFS[16'h202F] = 8'h02;
DFS[16'h2030] = 8'h0D;
DFS[16'h2031] = 8'h20;
DFS[16'h2032] = 8'h7B;
DFS[16'h2033] = 8'hA1;
DFS[16'h2034] = 8'h68;
DFS[16'h2035] = 8'h85;
DFS[16'h2036] = 8'hB8;
DFS[16'h2037] = 8'h68;
DFS[16'h2038] = 8'h85;
DFS[16'h2039] = 8'hB9;
DFS[16'h203A] = 8'h20;
DFS[16'h203B] = 8'h0F;
DFS[16'h203C] = 8'hA0;
DFS[16'h203D] = 8'hA5;
DFS[16'h203E] = 8'hB0;
DFS[16'h203F] = 8'h20;
DFS[16'h2040] = 8'h69;
DFS[16'h2041] = 8'hA0;
DFS[16'h2042] = 8'hA5;
DFS[16'h2043] = 8'hB1;
DFS[16'h2044] = 8'hF0;
DFS[16'h2045] = 8'h1B;
DFS[16'h2046] = 8'hA9;
DFS[16'h2047] = 8'h2F;
DFS[16'h2048] = 8'h99;
DFS[16'h2049] = 8'h00;
DFS[16'h204A] = 8'h01;
DFS[16'h204B] = 8'hC8;
DFS[16'h204C] = 8'hAE;
DFS[16'h204D] = 8'h41;
DFS[16'h204E] = 8'h0D;
DFS[16'h204F] = 8'hBD;
DFS[16'h2050] = 8'h44;
DFS[16'h2051] = 8'h0D;
DFS[16'h2052] = 8'h20;
DFS[16'h2053] = 8'h69;
DFS[16'h2054] = 8'hA0;
DFS[16'h2055] = 8'hBD;
DFS[16'h2056] = 8'h45;
DFS[16'h2057] = 8'h0D;
DFS[16'h2058] = 8'h20;
DFS[16'h2059] = 8'h69;
DFS[16'h205A] = 8'hA0;
DFS[16'h205B] = 8'hBD;
DFS[16'h205C] = 8'h46;
DFS[16'h205D] = 8'h0D;
DFS[16'h205E] = 8'h20;
DFS[16'h205F] = 8'h69;
DFS[16'h2060] = 8'hA0;
DFS[16'h2061] = 8'hA9;
DFS[16'h2062] = 8'h00;
DFS[16'h2063] = 8'h99;
DFS[16'h2064] = 8'h00;
DFS[16'h2065] = 8'h01;
DFS[16'h2066] = 8'h4C;
DFS[16'h2067] = 8'h00;
DFS[16'h2068] = 8'h01;
DFS[16'h2069] = 8'h48;
DFS[16'h206A] = 8'h4A;
DFS[16'h206B] = 8'h4A;
DFS[16'h206C] = 8'h4A;
DFS[16'h206D] = 8'h4A;
DFS[16'h206E] = 8'h20;
DFS[16'h206F] = 8'h74;
DFS[16'h2070] = 8'hA0;
DFS[16'h2071] = 8'h68;
DFS[16'h2072] = 8'h29;
DFS[16'h2073] = 8'h0F;
DFS[16'h2074] = 8'h18;
DFS[16'h2075] = 8'h69;
DFS[16'h2076] = 8'h30;
DFS[16'h2077] = 8'hC9;
DFS[16'h2078] = 8'h3A;
DFS[16'h2079] = 8'h90;
DFS[16'h207A] = 8'h02;
DFS[16'h207B] = 8'h69;
DFS[16'h207C] = 8'h06;
DFS[16'h207D] = 8'h99;
DFS[16'h207E] = 8'h00;
DFS[16'h207F] = 8'h01;
DFS[16'h2080] = 8'hC8;
DFS[16'h2081] = 8'h60;
DFS[16'h2082] = 8'h20;
DFS[16'h2083] = 8'h00;
DFS[16'h2084] = 8'hA0;
DFS[16'h2085] = 8'h11;
DFS[16'h2086] = 8'h45;
DFS[16'h2087] = 8'h73;
DFS[16'h2088] = 8'h63;
DFS[16'h2089] = 8'h61;
DFS[16'h208A] = 8'h70;
DFS[16'h208B] = 8'h65;
DFS[16'h208C] = 8'h00;
DFS[16'h208D] = 8'h48;
DFS[16'h208E] = 8'hA9;
DFS[16'h208F] = 8'hFF;
DFS[16'h2090] = 8'h8D;
DFS[16'h2091] = 8'h74;
DFS[16'h2092] = 8'h10;
DFS[16'h2093] = 8'h8D;
DFS[16'h2094] = 8'h75;
DFS[16'h2095] = 8'h10;
DFS[16'h2096] = 8'h68;
DFS[16'h2097] = 8'h60;
DFS[16'h2098] = 8'h48;
DFS[16'h2099] = 8'hA5;
DFS[16'h209A] = 8'hBE;
DFS[16'h209B] = 8'h8D;
DFS[16'h209C] = 8'h72;
DFS[16'h209D] = 8'h10;
DFS[16'h209E] = 8'hA5;
DFS[16'h209F] = 8'hBF;
DFS[16'h20A0] = 8'h8D;
DFS[16'h20A1] = 8'h73;
DFS[16'h20A2] = 8'h10;
DFS[16'h20A3] = 8'hAD;
DFS[16'h20A4] = 8'h74;
DFS[16'h20A5] = 8'h10;
DFS[16'h20A6] = 8'h2D;
DFS[16'h20A7] = 8'h75;
DFS[16'h20A8] = 8'h10;
DFS[16'h20A9] = 8'h0D;
DFS[16'h20AA] = 8'hD7;
DFS[16'h20AB] = 8'h10;
DFS[16'h20AC] = 8'h49;
DFS[16'h20AD] = 8'hFF;
DFS[16'h20AE] = 8'h8D;
DFS[16'h20AF] = 8'hD6;
DFS[16'h20B0] = 8'h10;
DFS[16'h20B1] = 8'h38;
DFS[16'h20B2] = 8'hF0;
DFS[16'h20B3] = 8'h0D;
DFS[16'h20B4] = 8'h20;
DFS[16'h20B5] = 8'hC3;
DFS[16'h20B6] = 8'hA0;
DFS[16'h20B7] = 8'hA2;
DFS[16'h20B8] = 8'h72;
DFS[16'h20B9] = 8'hA0;
DFS[16'h20BA] = 8'h10;
DFS[16'h20BB] = 8'h68;
DFS[16'h20BC] = 8'h48;
DFS[16'h20BD] = 8'h20;
DFS[16'h20BE] = 8'h06;
DFS[16'h20BF] = 8'h04;
DFS[16'h20C0] = 8'h18;
DFS[16'h20C1] = 8'h68;
DFS[16'h20C2] = 8'h60;
DFS[16'h20C3] = 8'h48;
DFS[16'h20C4] = 8'hA9;
DFS[16'h20C5] = 8'hC1;
DFS[16'h20C6] = 8'h20;
DFS[16'h20C7] = 8'h06;
DFS[16'h20C8] = 8'h04;
DFS[16'h20C9] = 8'h90;
DFS[16'h20CA] = 8'hF9;
DFS[16'h20CB] = 8'h68;
DFS[16'h20CC] = 8'h60;
DFS[16'h20CD] = 8'hAD;
DFS[16'h20CE] = 8'hD6;
DFS[16'h20CF] = 8'h10;
DFS[16'h20D0] = 8'hF0;
DFS[16'h20D1] = 8'h05;
DFS[16'h20D2] = 8'hA9;
DFS[16'h20D3] = 8'h81;
DFS[16'h20D4] = 8'h20;
DFS[16'h20D5] = 8'h06;
DFS[16'h20D6] = 8'h04;
DFS[16'h20D7] = 8'h60;
DFS[16'h20D8] = 8'h9D;
DFS[16'h20D9] = 8'h05;
DFS[16'h20DA] = 8'h01;
DFS[16'h20DB] = 8'h20;
DFS[16'h20DC] = 8'hE4;
DFS[16'h20DD] = 8'h95;
DFS[16'h20DE] = 8'h08;
DFS[16'h20DF] = 8'hAD;
DFS[16'h20E0] = 8'h81;
DFS[16'h20E1] = 8'h10;
DFS[16'h20E2] = 8'hF0;
DFS[16'h20E3] = 8'h05;
DFS[16'h20E4] = 8'hA9;
DFS[16'h20E5] = 8'h81;
DFS[16'h20E6] = 8'h20;
DFS[16'h20E7] = 8'h06;
DFS[16'h20E8] = 8'h04;
DFS[16'h20E9] = 8'h28;
DFS[16'h20EA] = 8'h60;
DFS[16'h20EB] = 8'hF0;
DFS[16'h20EC] = 8'h06;
DFS[16'h20ED] = 8'h20;
DFS[16'h20EE] = 8'hC3;
DFS[16'h20EF] = 8'hA0;
DFS[16'h20F0] = 8'h18;
DFS[16'h20F1] = 8'hA9;
DFS[16'h20F2] = 8'hFF;
DFS[16'h20F3] = 8'h4C;
DFS[16'h20F4] = 8'h17;
DFS[16'h20F5] = 8'h96;
DFS[16'h20F6] = 8'hC9;
DFS[16'h20F7] = 8'hFE;
DFS[16'h20F8] = 8'h90;
DFS[16'h20F9] = 8'h5A;
DFS[16'h20FA] = 8'hD0;
DFS[16'h20FB] = 8'h1B;
DFS[16'h20FC] = 8'hC0;
DFS[16'h20FD] = 8'h00;
DFS[16'h20FE] = 8'hF0;
DFS[16'h20FF] = 8'h54;
DFS[16'h2100] = 8'hA2;
DFS[16'h2101] = 8'h06;
DFS[16'h2102] = 8'hA9;
DFS[16'h2103] = 8'h14;
DFS[16'h2104] = 8'h20;
DFS[16'h2105] = 8'hF4;
DFS[16'h2106] = 8'hFF;
DFS[16'h2107] = 8'h2C;
DFS[16'h2108] = 8'hE0;
DFS[16'h2109] = 8'hFE;
DFS[16'h210A] = 8'h10;
DFS[16'h210B] = 8'hFB;
DFS[16'h210C] = 8'hAD;
DFS[16'h210D] = 8'hE1;
DFS[16'h210E] = 8'hFE;
DFS[16'h210F] = 8'hF0;
DFS[16'h2110] = 8'h41;
DFS[16'h2111] = 8'h20;
DFS[16'h2112] = 8'hEE;
DFS[16'h2113] = 8'hFF;
DFS[16'h2114] = 8'h4C;
DFS[16'h2115] = 8'h07;
DFS[16'h2116] = 8'hA1;
DFS[16'h2117] = 8'hA9;
DFS[16'h2118] = 8'hAD;
DFS[16'h2119] = 8'h8D;
DFS[16'h211A] = 8'h20;
DFS[16'h211B] = 8'h02;
DFS[16'h211C] = 8'hA9;
DFS[16'h211D] = 8'h06;
DFS[16'h211E] = 8'h8D;
DFS[16'h211F] = 8'h21;
DFS[16'h2120] = 8'h02;
DFS[16'h2121] = 8'hA9;
DFS[16'h2122] = 8'h16;
DFS[16'h2123] = 8'h8D;
DFS[16'h2124] = 8'h02;
DFS[16'h2125] = 8'h02;
DFS[16'h2126] = 8'hA0;
DFS[16'h2127] = 8'h00;
DFS[16'h2128] = 8'h8C;
DFS[16'h2129] = 8'h03;
DFS[16'h212A] = 8'h02;
DFS[16'h212B] = 8'hA9;
DFS[16'h212C] = 8'h8E;
DFS[16'h212D] = 8'h8D;
DFS[16'h212E] = 8'hE0;
DFS[16'h212F] = 8'hFE;
DFS[16'h2130] = 8'hB9;
DFS[16'h2131] = 8'h03;
DFS[16'h2132] = 8'h8B;
DFS[16'h2133] = 8'h99;
DFS[16'h2134] = 8'h00;
DFS[16'h2135] = 8'h04;
DFS[16'h2136] = 8'hB9;
DFS[16'h2137] = 8'h03;
DFS[16'h2138] = 8'h8C;
DFS[16'h2139] = 8'h99;
DFS[16'h213A] = 8'h00;
DFS[16'h213B] = 8'h05;
DFS[16'h213C] = 8'hB9;
DFS[16'h213D] = 8'h03;
DFS[16'h213E] = 8'h8D;
DFS[16'h213F] = 8'h99;
DFS[16'h2140] = 8'h00;
DFS[16'h2141] = 8'h06;
DFS[16'h2142] = 8'h88;
DFS[16'h2143] = 8'hD0;
DFS[16'h2144] = 8'hEB;
DFS[16'h2145] = 8'h20;
DFS[16'h2146] = 8'h21;
DFS[16'h2147] = 8'h04;
DFS[16'h2148] = 8'hA2;
DFS[16'h2149] = 8'h40;
DFS[16'h214A] = 8'hBD;
DFS[16'h214B] = 8'hC2;
DFS[16'h214C] = 8'h8A;
DFS[16'h214D] = 8'h95;
DFS[16'h214E] = 8'h16;
DFS[16'h214F] = 8'hCA;
DFS[16'h2150] = 8'h10;
DFS[16'h2151] = 8'hF8;
DFS[16'h2152] = 8'hA9;
DFS[16'h2153] = 8'h00;
DFS[16'h2154] = 8'h60;
DFS[16'h2155] = 8'hA9;
DFS[16'h2156] = 8'hFF;
DFS[16'h2157] = 8'h8D;
DFS[16'h2158] = 8'h52;
DFS[16'h2159] = 8'h0D;
DFS[16'h215A] = 8'h48;
DFS[16'h215B] = 8'h4C;
DFS[16'h215C] = 8'h3B;
DFS[16'h215D] = 8'h93;
DFS[16'h215E] = 8'hB9;
DFS[16'h215F] = 8'h14;
DFS[16'h2160] = 8'h11;
DFS[16'h2161] = 8'h99;
DFS[16'h2162] = 8'h10;
DFS[16'h2163] = 8'h11;
DFS[16'h2164] = 8'hB9;
DFS[16'h2165] = 8'h15;
DFS[16'h2166] = 8'h11;
DFS[16'h2167] = 8'h99;
DFS[16'h2168] = 8'h11;
DFS[16'h2169] = 8'h11;
DFS[16'h216A] = 8'hB9;
DFS[16'h216B] = 8'h16;
DFS[16'h216C] = 8'h11;
DFS[16'h216D] = 8'h99;
DFS[16'h216E] = 8'h12;
DFS[16'h216F] = 8'h11;
DFS[16'h2170] = 8'h60;
DFS[16'h2171] = 8'hA2;
DFS[16'h2172] = 8'h06;
DFS[16'h2173] = 8'h8E;
DFS[16'h2174] = 8'h40;
DFS[16'h2175] = 8'hFE;
DFS[16'h2176] = 8'hE8;
DFS[16'h2177] = 8'h8E;
DFS[16'h2178] = 8'h40;
DFS[16'h2179] = 8'hFE;
DFS[16'h217A] = 8'h60;
DFS[16'h217B] = 8'hA9;
DFS[16'h217C] = 8'h76;
DFS[16'h217D] = 8'h4C;
DFS[16'h217E] = 8'hF4;
DFS[16'h217F] = 8'hFF;
DFS[16'h2180] = 8'hA2;
DFS[16'h2181] = 8'h01;
DFS[16'h2182] = 8'hA9;
DFS[16'h2183] = 8'h03;
DFS[16'h2184] = 8'h8E;
DFS[16'h2185] = 8'h60;
DFS[16'h2186] = 8'hFE;
DFS[16'h2187] = 8'h8D;
DFS[16'h2188] = 8'h60;
DFS[16'h2189] = 8'hFE;
DFS[16'h218A] = 8'h8E;
DFS[16'h218B] = 8'h60;
DFS[16'h218C] = 8'hFE;
DFS[16'h218D] = 8'h8D;
DFS[16'h218E] = 8'h60;
DFS[16'h218F] = 8'hFE;
DFS[16'h2190] = 8'h8E;
DFS[16'h2191] = 8'h60;
DFS[16'h2192] = 8'hFE;
DFS[16'h2193] = 8'h8D;
DFS[16'h2194] = 8'h60;
DFS[16'h2195] = 8'hFE;
DFS[16'h2196] = 8'h8E;
DFS[16'h2197] = 8'h60;
DFS[16'h2198] = 8'hFE;
DFS[16'h2199] = 8'h8D;
DFS[16'h219A] = 8'h60;
DFS[16'h219B] = 8'hFE;
DFS[16'h219C] = 8'h8E;
DFS[16'h219D] = 8'h60;
DFS[16'h219E] = 8'hFE;
DFS[16'h219F] = 8'h8D;
DFS[16'h21A0] = 8'h60;
DFS[16'h21A1] = 8'hFE;
DFS[16'h21A2] = 8'h8E;
DFS[16'h21A3] = 8'h60;
DFS[16'h21A4] = 8'hFE;
DFS[16'h21A5] = 8'h8D;
DFS[16'h21A6] = 8'h60;
DFS[16'h21A7] = 8'hFE;
DFS[16'h21A8] = 8'h8E;
DFS[16'h21A9] = 8'h60;
DFS[16'h21AA] = 8'hFE;
DFS[16'h21AB] = 8'h8D;
DFS[16'h21AC] = 8'h60;
DFS[16'h21AD] = 8'hFE;
DFS[16'h21AE] = 8'h8E;
DFS[16'h21AF] = 8'h60;
DFS[16'h21B0] = 8'hFE;
DFS[16'h21B1] = 8'h8D;
DFS[16'h21B2] = 8'h60;
DFS[16'h21B3] = 8'hFE;
DFS[16'h21B4] = 8'hAD;
DFS[16'h21B5] = 8'h6A;
DFS[16'h21B6] = 8'hFE;
DFS[16'h21B7] = 8'h60;
DFS[16'h21B8] = 8'h0A;
DFS[16'h21B9] = 8'h2A;
DFS[16'h21BA] = 8'h8D;
DFS[16'h21BB] = 8'h60;
DFS[16'h21BC] = 8'hFE;
DFS[16'h21BD] = 8'h09;
DFS[16'h21BE] = 8'h02;
DFS[16'h21BF] = 8'h8D;
DFS[16'h21C0] = 8'h60;
DFS[16'h21C1] = 8'hFE;
DFS[16'h21C2] = 8'h2A;
DFS[16'h21C3] = 8'h29;
DFS[16'h21C4] = 8'hFD;
DFS[16'h21C5] = 8'h8D;
DFS[16'h21C6] = 8'h60;
DFS[16'h21C7] = 8'hFE;
DFS[16'h21C8] = 8'h09;
DFS[16'h21C9] = 8'h02;
DFS[16'h21CA] = 8'h8D;
DFS[16'h21CB] = 8'h60;
DFS[16'h21CC] = 8'hFE;
DFS[16'h21CD] = 8'h2A;
DFS[16'h21CE] = 8'h29;
DFS[16'h21CF] = 8'hFD;
DFS[16'h21D0] = 8'h8D;
DFS[16'h21D1] = 8'h60;
DFS[16'h21D2] = 8'hFE;
DFS[16'h21D3] = 8'h09;
DFS[16'h21D4] = 8'h02;
DFS[16'h21D5] = 8'h8D;
DFS[16'h21D6] = 8'h60;
DFS[16'h21D7] = 8'hFE;
DFS[16'h21D8] = 8'h2A;
DFS[16'h21D9] = 8'h29;
DFS[16'h21DA] = 8'hFD;
DFS[16'h21DB] = 8'h8D;
DFS[16'h21DC] = 8'h60;
DFS[16'h21DD] = 8'hFE;
DFS[16'h21DE] = 8'h09;
DFS[16'h21DF] = 8'h02;
DFS[16'h21E0] = 8'h8D;
DFS[16'h21E1] = 8'h60;
DFS[16'h21E2] = 8'hFE;
DFS[16'h21E3] = 8'h2A;
DFS[16'h21E4] = 8'h29;
DFS[16'h21E5] = 8'hFD;
DFS[16'h21E6] = 8'h8D;
DFS[16'h21E7] = 8'h60;
DFS[16'h21E8] = 8'hFE;
DFS[16'h21E9] = 8'h09;
DFS[16'h21EA] = 8'h02;
DFS[16'h21EB] = 8'h8D;
DFS[16'h21EC] = 8'h60;
DFS[16'h21ED] = 8'hFE;
DFS[16'h21EE] = 8'h2A;
DFS[16'h21EF] = 8'h29;
DFS[16'h21F0] = 8'hFD;
DFS[16'h21F1] = 8'h8D;
DFS[16'h21F2] = 8'h60;
DFS[16'h21F3] = 8'hFE;
DFS[16'h21F4] = 8'h09;
DFS[16'h21F5] = 8'h02;
DFS[16'h21F6] = 8'h8D;
DFS[16'h21F7] = 8'h60;
DFS[16'h21F8] = 8'hFE;
DFS[16'h21F9] = 8'h2A;
DFS[16'h21FA] = 8'h29;
DFS[16'h21FB] = 8'hFD;
DFS[16'h21FC] = 8'h8D;
DFS[16'h21FD] = 8'h60;
DFS[16'h21FE] = 8'hFE;
DFS[16'h21FF] = 8'h09;
DFS[16'h2200] = 8'h02;
DFS[16'h2201] = 8'h8D;
DFS[16'h2202] = 8'h60;
DFS[16'h2203] = 8'hFE;
DFS[16'h2204] = 8'h2A;
DFS[16'h2205] = 8'h29;
DFS[16'h2206] = 8'hFD;
DFS[16'h2207] = 8'h8D;
DFS[16'h2208] = 8'h60;
DFS[16'h2209] = 8'hFE;
DFS[16'h220A] = 8'h09;
DFS[16'h220B] = 8'h02;
DFS[16'h220C] = 8'h8D;
DFS[16'h220D] = 8'h60;
DFS[16'h220E] = 8'hFE;
DFS[16'h220F] = 8'h60;
DFS[16'h2210] = 8'h2C;
DFS[16'h2211] = 8'h40;
DFS[16'h2212] = 8'h0D;
DFS[16'h2213] = 8'h30;
DFS[16'h2214] = 8'h38;
DFS[16'h2215] = 8'hA2;
DFS[16'h2216] = 8'h01;
DFS[16'h2217] = 8'hA9;
DFS[16'h2218] = 8'h03;
DFS[16'h2219] = 8'h8E;
DFS[16'h221A] = 8'h60;
DFS[16'h221B] = 8'hFE;
DFS[16'h221C] = 8'h8D;
DFS[16'h221D] = 8'h60;
DFS[16'h221E] = 8'hFE;
DFS[16'h221F] = 8'h8E;
DFS[16'h2220] = 8'h60;
DFS[16'h2221] = 8'hFE;
DFS[16'h2222] = 8'h8D;
DFS[16'h2223] = 8'h60;
DFS[16'h2224] = 8'hFE;
DFS[16'h2225] = 8'h8E;
DFS[16'h2226] = 8'h60;
DFS[16'h2227] = 8'hFE;
DFS[16'h2228] = 8'h8D;
DFS[16'h2229] = 8'h60;
DFS[16'h222A] = 8'hFE;
DFS[16'h222B] = 8'h8E;
DFS[16'h222C] = 8'h60;
DFS[16'h222D] = 8'hFE;
DFS[16'h222E] = 8'h8D;
DFS[16'h222F] = 8'h60;
DFS[16'h2230] = 8'hFE;
DFS[16'h2231] = 8'h8E;
DFS[16'h2232] = 8'h60;
DFS[16'h2233] = 8'hFE;
DFS[16'h2234] = 8'h8D;
DFS[16'h2235] = 8'h60;
DFS[16'h2236] = 8'hFE;
DFS[16'h2237] = 8'h8E;
DFS[16'h2238] = 8'h60;
DFS[16'h2239] = 8'hFE;
DFS[16'h223A] = 8'h8D;
DFS[16'h223B] = 8'h60;
DFS[16'h223C] = 8'hFE;
DFS[16'h223D] = 8'h8E;
DFS[16'h223E] = 8'h60;
DFS[16'h223F] = 8'hFE;
DFS[16'h2240] = 8'h8D;
DFS[16'h2241] = 8'h60;
DFS[16'h2242] = 8'hFE;
DFS[16'h2243] = 8'h8E;
DFS[16'h2244] = 8'h60;
DFS[16'h2245] = 8'hFE;
DFS[16'h2246] = 8'h8D;
DFS[16'h2247] = 8'h60;
DFS[16'h2248] = 8'hFE;
DFS[16'h2249] = 8'h88;
DFS[16'h224A] = 8'hD0;
DFS[16'h224B] = 8'hCD;
DFS[16'h224C] = 8'h60;
DFS[16'h224D] = 8'hA9;
DFS[16'h224E] = 8'hFF;
DFS[16'h224F] = 8'h8D;
DFS[16'h2250] = 8'h18;
DFS[16'h2251] = 8'hFE;
DFS[16'h2252] = 8'hEA;
DFS[16'h2253] = 8'hEA;
DFS[16'h2254] = 8'hEA;
DFS[16'h2255] = 8'h88;
DFS[16'h2256] = 8'hD0;
DFS[16'h2257] = 8'hF7;
DFS[16'h2258] = 8'h60;
DFS[16'h2259] = 8'h2C;
DFS[16'h225A] = 8'h40;
DFS[16'h225B] = 8'h0D;
DFS[16'h225C] = 8'h30;
DFS[16'h225D] = 8'h36;
DFS[16'h225E] = 8'h8E;
DFS[16'h225F] = 8'h41;
DFS[16'h2260] = 8'h0D;
DFS[16'h2261] = 8'hA0;
DFS[16'h2262] = 8'h07;
DFS[16'h2263] = 8'hBD;
DFS[16'h2264] = 8'h42;
DFS[16'h2265] = 8'h0D;
DFS[16'h2266] = 8'h20;
DFS[16'h2267] = 8'hB8;
DFS[16'h2268] = 8'hA1;
DFS[16'h2269] = 8'hE8;
DFS[16'h226A] = 8'h88;
DFS[16'h226B] = 8'hD0;
DFS[16'h226C] = 8'hF6;
DFS[16'h226D] = 8'h20;
DFS[16'h226E] = 8'h73;
DFS[16'h226F] = 8'hA2;
DFS[16'h2270] = 8'h4C;
DFS[16'h2271] = 8'h8A;
DFS[16'h2272] = 8'hA1;
DFS[16'h2273] = 8'hA9;
DFS[16'h2274] = 8'h01;
DFS[16'h2275] = 8'hA2;
DFS[16'h2276] = 8'h03;
DFS[16'h2277] = 8'hA0;
DFS[16'h2278] = 8'h00;
DFS[16'h2279] = 8'h88;
DFS[16'h227A] = 8'hF0;
DFS[16'h227B] = 8'h12;
DFS[16'h227C] = 8'h8D;
DFS[16'h227D] = 8'h60;
DFS[16'h227E] = 8'hFE;
DFS[16'h227F] = 8'h8E;
DFS[16'h2280] = 8'h60;
DFS[16'h2281] = 8'hFE;
DFS[16'h2282] = 8'hAD;
DFS[16'h2283] = 8'h6A;
DFS[16'h2284] = 8'hFE;
DFS[16'h2285] = 8'h29;
DFS[16'h2286] = 8'h01;
DFS[16'h2287] = 8'hD0;
DFS[16'h2288] = 8'hF0;
DFS[16'h2289] = 8'hA2;
DFS[16'h228A] = 8'h01;
DFS[16'h228B] = 8'hA9;
DFS[16'h228C] = 8'h03;
DFS[16'h228D] = 8'h60;
DFS[16'h228E] = 8'hAD;
DFS[16'h228F] = 8'h6A;
DFS[16'h2290] = 8'hFE;
DFS[16'h2291] = 8'hC9;
DFS[16'h2292] = 8'h00;
DFS[16'h2293] = 8'h60;
DFS[16'h2294] = 8'h8E;
DFS[16'h2295] = 8'h41;
DFS[16'h2296] = 8'h0D;
DFS[16'h2297] = 8'hA0;
DFS[16'h2298] = 8'h08;
DFS[16'h2299] = 8'hBD;
DFS[16'h229A] = 8'h42;
DFS[16'h229B] = 8'h0D;
DFS[16'h229C] = 8'h8D;
DFS[16'h229D] = 8'h18;
DFS[16'h229E] = 8'hFE;
DFS[16'h229F] = 8'hEA;
DFS[16'h22A0] = 8'hEA;
DFS[16'h22A1] = 8'hE8;
DFS[16'h22A2] = 8'h88;
DFS[16'h22A3] = 8'hD0;
DFS[16'h22A4] = 8'hF4;
DFS[16'h22A5] = 8'h8D;
DFS[16'h22A6] = 8'h18;
DFS[16'h22A7] = 8'hFE;
DFS[16'h22A8] = 8'h20;
DFS[16'h22A9] = 8'h58;
DFS[16'h22AA] = 8'hA2;
DFS[16'h22AB] = 8'hAD;
DFS[16'h22AC] = 8'h18;
DFS[16'h22AD] = 8'hFE;
DFS[16'h22AE] = 8'h10;
DFS[16'h22AF] = 8'hE3;
DFS[16'h22B0] = 8'h88;
DFS[16'h22B1] = 8'hD0;
DFS[16'h22B2] = 8'hF5;
DFS[16'h22B3] = 8'h4C;
DFS[16'h22B4] = 8'h91;
DFS[16'h22B5] = 8'hA2;
DFS[16'h22B6] = 8'h2C;
DFS[16'h22B7] = 8'h40;
DFS[16'h22B8] = 8'h0D;
DFS[16'h22B9] = 8'h30;
DFS[16'h22BA] = 8'h0A;
DFS[16'h22BB] = 8'hA2;
DFS[16'h22BC] = 8'h01;
DFS[16'h22BD] = 8'h20;
DFS[16'h22BE] = 8'h82;
DFS[16'h22BF] = 8'hA1;
DFS[16'h22C0] = 8'hC9;
DFS[16'h22C1] = 8'hFE;
DFS[16'h22C2] = 8'hD0;
DFS[16'h22C3] = 8'hF9;
DFS[16'h22C4] = 8'h60;
DFS[16'h22C5] = 8'hA2;
DFS[16'h22C6] = 8'hFF;
DFS[16'h22C7] = 8'h8E;
DFS[16'h22C8] = 8'h18;
DFS[16'h22C9] = 8'hFE;
DFS[16'h22CA] = 8'h20;
DFS[16'h22CB] = 8'h58;
DFS[16'h22CC] = 8'hA2;
DFS[16'h22CD] = 8'hAD;
DFS[16'h22CE] = 8'h18;
DFS[16'h22CF] = 8'hFE;
DFS[16'h22D0] = 8'hC9;
DFS[16'h22D1] = 8'hFE;
DFS[16'h22D2] = 8'hD0;
DFS[16'h22D3] = 8'hF3;
DFS[16'h22D4] = 8'h60;
DFS[16'h22D5] = 8'h2C;
DFS[16'h22D6] = 8'h40;
DFS[16'h22D7] = 8'h0D;
DFS[16'h22D8] = 8'h30;
DFS[16'h22D9] = 8'h15;
DFS[16'h22DA] = 8'hA2;
DFS[16'h22DB] = 8'h01;
DFS[16'h22DC] = 8'hAC;
DFS[16'h22DD] = 8'hD6;
DFS[16'h22DE] = 8'h10;
DFS[16'h22DF] = 8'hD0;
DFS[16'h22E0] = 8'h09;
DFS[16'h22E1] = 8'h20;
DFS[16'h22E2] = 8'h82;
DFS[16'h22E3] = 8'hA1;
DFS[16'h22E4] = 8'h91;
DFS[16'h22E5] = 8'hA0;
DFS[16'h22E6] = 8'hC8;
DFS[16'h22E7] = 8'hD0;
DFS[16'h22E8] = 8'hF8;
DFS[16'h22E9] = 8'h60;
DFS[16'h22EA] = 8'hA0;
DFS[16'h22EB] = 8'h00;
DFS[16'h22EC] = 8'h4C;
DFS[16'h22ED] = 8'h2D;
DFS[16'h22EE] = 8'hA3;
DFS[16'h22EF] = 8'hA2;
DFS[16'h22F0] = 8'hFF;
DFS[16'h22F1] = 8'h8E;
DFS[16'h22F2] = 8'h18;
DFS[16'h22F3] = 8'hFE;
DFS[16'h22F4] = 8'hAC;
DFS[16'h22F5] = 8'hD6;
DFS[16'h22F6] = 8'h10;
DFS[16'h22F7] = 8'hD0;
DFS[16'h22F8] = 8'h16;
DFS[16'h22F9] = 8'hEA;
DFS[16'h22FA] = 8'hEA;
DFS[16'h22FB] = 8'hEA;
DFS[16'h22FC] = 8'hAD;
DFS[16'h22FD] = 8'h18;
DFS[16'h22FE] = 8'hFE;
DFS[16'h22FF] = 8'h8E;
DFS[16'h2300] = 8'h18;
DFS[16'h2301] = 8'hFE;
DFS[16'h2302] = 8'h91;
DFS[16'h2303] = 8'hA0;
DFS[16'h2304] = 8'hC8;
DFS[16'h2305] = 8'hC0;
DFS[16'h2306] = 8'hFF;
DFS[16'h2307] = 8'hD0;
DFS[16'h2308] = 8'hF3;
DFS[16'h2309] = 8'hAD;
DFS[16'h230A] = 8'h18;
DFS[16'h230B] = 8'hFE;
DFS[16'h230C] = 8'h91;
DFS[16'h230D] = 8'hA0;
DFS[16'h230E] = 8'h60;
DFS[16'h230F] = 8'hA0;
DFS[16'h2310] = 8'h00;
DFS[16'h2311] = 8'h4C;
DFS[16'h2312] = 8'h5A;
DFS[16'h2313] = 8'hA3;
DFS[16'h2314] = 8'h2C;
DFS[16'h2315] = 8'h40;
DFS[16'h2316] = 8'h0D;
DFS[16'h2317] = 8'h30;
DFS[16'h2318] = 8'h1E;
DFS[16'h2319] = 8'hA2;
DFS[16'h231A] = 8'h01;
DFS[16'h231B] = 8'hAC;
DFS[16'h231C] = 8'hD6;
DFS[16'h231D] = 8'h10;
DFS[16'h231E] = 8'hD0;
DFS[16'h231F] = 8'h0B;
DFS[16'h2320] = 8'h20;
DFS[16'h2321] = 8'h82;
DFS[16'h2322] = 8'hA1;
DFS[16'h2323] = 8'h91;
DFS[16'h2324] = 8'hA0;
DFS[16'h2325] = 8'hC8;
DFS[16'h2326] = 8'hC6;
DFS[16'h2327] = 8'hA7;
DFS[16'h2328] = 8'hD0;
DFS[16'h2329] = 8'hF6;
DFS[16'h232A] = 8'h60;
DFS[16'h232B] = 8'hA4;
DFS[16'h232C] = 8'hA7;
DFS[16'h232D] = 8'h20;
DFS[16'h232E] = 8'h82;
DFS[16'h232F] = 8'hA1;
DFS[16'h2330] = 8'h8D;
DFS[16'h2331] = 8'hE5;
DFS[16'h2332] = 8'hFE;
DFS[16'h2333] = 8'h88;
DFS[16'h2334] = 8'hD0;
DFS[16'h2335] = 8'hF7;
DFS[16'h2336] = 8'h60;
DFS[16'h2337] = 8'hA2;
DFS[16'h2338] = 8'hFF;
DFS[16'h2339] = 8'h8E;
DFS[16'h233A] = 8'h18;
DFS[16'h233B] = 8'hFE;
DFS[16'h233C] = 8'hAC;
DFS[16'h233D] = 8'hD6;
DFS[16'h233E] = 8'h10;
DFS[16'h233F] = 8'hD0;
DFS[16'h2340] = 8'h17;
DFS[16'h2341] = 8'hC6;
DFS[16'h2342] = 8'hA7;
DFS[16'h2343] = 8'hF0;
DFS[16'h2344] = 8'h0D;
DFS[16'h2345] = 8'hAD;
DFS[16'h2346] = 8'h18;
DFS[16'h2347] = 8'hFE;
DFS[16'h2348] = 8'h8E;
DFS[16'h2349] = 8'h18;
DFS[16'h234A] = 8'hFE;
DFS[16'h234B] = 8'h91;
DFS[16'h234C] = 8'hA0;
DFS[16'h234D] = 8'hC8;
DFS[16'h234E] = 8'hC6;
DFS[16'h234F] = 8'hA7;
DFS[16'h2350] = 8'hD0;
DFS[16'h2351] = 8'hF3;
DFS[16'h2352] = 8'hAD;
DFS[16'h2353] = 8'h18;
DFS[16'h2354] = 8'hFE;
DFS[16'h2355] = 8'h91;
DFS[16'h2356] = 8'hA0;
DFS[16'h2357] = 8'h60;
DFS[16'h2358] = 8'hA4;
DFS[16'h2359] = 8'hA7;
DFS[16'h235A] = 8'h88;
DFS[16'h235B] = 8'hF0;
DFS[16'h235C] = 8'h1A;
DFS[16'h235D] = 8'hEA;
DFS[16'h235E] = 8'hAD;
DFS[16'h235F] = 8'h18;
DFS[16'h2360] = 8'hFE;
DFS[16'h2361] = 8'h8E;
DFS[16'h2362] = 8'h18;
DFS[16'h2363] = 8'hFE;
DFS[16'h2364] = 8'h8D;
DFS[16'h2365] = 8'hE5;
DFS[16'h2366] = 8'hFE;
DFS[16'h2367] = 8'h20;
DFS[16'h2368] = 8'h58;
DFS[16'h2369] = 8'hA2;
DFS[16'h236A] = 8'h20;
DFS[16'h236B] = 8'h58;
DFS[16'h236C] = 8'hA2;
DFS[16'h236D] = 8'hEA;
DFS[16'h236E] = 8'hEA;
DFS[16'h236F] = 8'hEA;
DFS[16'h2370] = 8'h88;
DFS[16'h2371] = 8'hD0;
DFS[16'h2372] = 8'hEA;
DFS[16'h2373] = 8'hEA;
DFS[16'h2374] = 8'hEA;
DFS[16'h2375] = 8'hEA;
DFS[16'h2376] = 8'hEA;
DFS[16'h2377] = 8'hAD;
DFS[16'h2378] = 8'h18;
DFS[16'h2379] = 8'hFE;
DFS[16'h237A] = 8'h8D;
DFS[16'h237B] = 8'hE5;
DFS[16'h237C] = 8'hFE;
DFS[16'h237D] = 8'h60;
DFS[16'h237E] = 8'h2C;
DFS[16'h237F] = 8'h40;
DFS[16'h2380] = 8'h0D;
DFS[16'h2381] = 8'h30;
DFS[16'h2382] = 8'h0E;
DFS[16'h2383] = 8'hA0;
DFS[16'h2384] = 8'h00;
DFS[16'h2385] = 8'hA2;
DFS[16'h2386] = 8'h01;
DFS[16'h2387] = 8'h20;
DFS[16'h2388] = 8'h82;
DFS[16'h2389] = 8'hA1;
DFS[16'h238A] = 8'h99;
DFS[16'h238B] = 8'h00;
DFS[16'h238C] = 8'h0E;
DFS[16'h238D] = 8'hC8;
DFS[16'h238E] = 8'hD0;
DFS[16'h238F] = 8'hF7;
DFS[16'h2390] = 8'h60;
DFS[16'h2391] = 8'hA0;
DFS[16'h2392] = 8'h00;
DFS[16'h2393] = 8'hA2;
DFS[16'h2394] = 8'hFF;
DFS[16'h2395] = 8'h8E;
DFS[16'h2396] = 8'h18;
DFS[16'h2397] = 8'hFE;
DFS[16'h2398] = 8'h20;
DFS[16'h2399] = 8'h58;
DFS[16'h239A] = 8'hA2;
DFS[16'h239B] = 8'hAD;
DFS[16'h239C] = 8'h18;
DFS[16'h239D] = 8'hFE;
DFS[16'h239E] = 8'h8E;
DFS[16'h239F] = 8'h18;
DFS[16'h23A0] = 8'hFE;
DFS[16'h23A1] = 8'h99;
DFS[16'h23A2] = 8'h00;
DFS[16'h23A3] = 8'h0E;
DFS[16'h23A4] = 8'hC8;
DFS[16'h23A5] = 8'hC0;
DFS[16'h23A6] = 8'hFF;
DFS[16'h23A7] = 8'hD0;
DFS[16'h23A8] = 8'hF2;
DFS[16'h23A9] = 8'hAD;
DFS[16'h23AA] = 8'h18;
DFS[16'h23AB] = 8'hFE;
DFS[16'h23AC] = 8'h99;
DFS[16'h23AD] = 8'h00;
DFS[16'h23AE] = 8'h0E;
DFS[16'h23AF] = 8'h60;
DFS[16'h23B0] = 8'h2C;
DFS[16'h23B1] = 8'h40;
DFS[16'h23B2] = 8'h0D;
DFS[16'h23B3] = 8'h30;
DFS[16'h23B4] = 8'h0A;
DFS[16'h23B5] = 8'hA0;
DFS[16'h23B6] = 8'h02;
DFS[16'h23B7] = 8'h20;
DFS[16'h23B8] = 8'h15;
DFS[16'h23B9] = 8'hA2;
DFS[16'h23BA] = 8'hA9;
DFS[16'h23BB] = 8'hFE;
DFS[16'h23BC] = 8'h4C;
DFS[16'h23BD] = 8'hB8;
DFS[16'h23BE] = 8'hA1;
DFS[16'h23BF] = 8'hA2;
DFS[16'h23C0] = 8'hFF;
DFS[16'h23C1] = 8'h8E;
DFS[16'h23C2] = 8'h18;
DFS[16'h23C3] = 8'hFE;
DFS[16'h23C4] = 8'h20;
DFS[16'h23C5] = 8'h58;
DFS[16'h23C6] = 8'hA2;
DFS[16'h23C7] = 8'h8E;
DFS[16'h23C8] = 8'h18;
DFS[16'h23C9] = 8'hFE;
DFS[16'h23CA] = 8'h20;
DFS[16'h23CB] = 8'h58;
DFS[16'h23CC] = 8'hA2;
DFS[16'h23CD] = 8'hCA;
DFS[16'h23CE] = 8'h8E;
DFS[16'h23CF] = 8'h18;
DFS[16'h23D0] = 8'hFE;
DFS[16'h23D1] = 8'h60;
DFS[16'h23D2] = 8'hA0;
DFS[16'h23D3] = 8'h02;
DFS[16'h23D4] = 8'h2C;
DFS[16'h23D5] = 8'h40;
DFS[16'h23D6] = 8'h0D;
DFS[16'h23D7] = 8'h30;
DFS[16'h23D8] = 8'h1A;
DFS[16'h23D9] = 8'h20;
DFS[16'h23DA] = 8'h15;
DFS[16'h23DB] = 8'hA2;
DFS[16'h23DC] = 8'h20;
DFS[16'h23DD] = 8'h73;
DFS[16'h23DE] = 8'hA2;
DFS[16'h23DF] = 8'h20;
DFS[16'h23E0] = 8'h9C;
DFS[16'h23E1] = 8'hA1;
DFS[16'h23E2] = 8'hA8;
DFS[16'h23E3] = 8'h29;
DFS[16'h23E4] = 8'h1F;
DFS[16'h23E5] = 8'hC9;
DFS[16'h23E6] = 8'h05;
DFS[16'h23E7] = 8'hD0;
DFS[16'h23E8] = 8'h2D;
DFS[16'h23E9] = 8'hA2;
DFS[16'h23EA] = 8'h01;
DFS[16'h23EB] = 8'h20;
DFS[16'h23EC] = 8'h82;
DFS[16'h23ED] = 8'hA1;
DFS[16'h23EE] = 8'hC9;
DFS[16'h23EF] = 8'hFF;
DFS[16'h23F0] = 8'hD0;
DFS[16'h23F1] = 8'hF9;
DFS[16'h23F2] = 8'h60;
DFS[16'h23F3] = 8'h20;
DFS[16'h23F4] = 8'h4D;
DFS[16'h23F5] = 8'hA2;
DFS[16'h23F6] = 8'hA2;
DFS[16'h23F7] = 8'hFF;
DFS[16'h23F8] = 8'h8E;
DFS[16'h23F9] = 8'h18;
DFS[16'h23FA] = 8'hFE;
DFS[16'h23FB] = 8'h20;
DFS[16'h23FC] = 8'h58;
DFS[16'h23FD] = 8'hA2;
DFS[16'h23FE] = 8'hAD;
DFS[16'h23FF] = 8'h18;
DFS[16'h2400] = 8'hFE;
DFS[16'h2401] = 8'hA8;
DFS[16'h2402] = 8'h29;
DFS[16'h2403] = 8'h1F;
DFS[16'h2404] = 8'hC9;
DFS[16'h2405] = 8'h05;
DFS[16'h2406] = 8'hD0;
DFS[16'h2407] = 8'h0E;
DFS[16'h2408] = 8'hA9;
DFS[16'h2409] = 8'hFF;
DFS[16'h240A] = 8'h8E;
DFS[16'h240B] = 8'h18;
DFS[16'h240C] = 8'hFE;
DFS[16'h240D] = 8'h20;
DFS[16'h240E] = 8'h58;
DFS[16'h240F] = 8'hA2;
DFS[16'h2410] = 8'hCD;
DFS[16'h2411] = 8'h18;
DFS[16'h2412] = 8'hFE;
DFS[16'h2413] = 8'hD0;
DFS[16'h2414] = 8'hF5;
DFS[16'h2415] = 8'h60;
DFS[16'h2416] = 8'h98;
DFS[16'h2417] = 8'h20;
DFS[16'h2418] = 8'h1F;
DFS[16'h2419] = 8'hA0;
DFS[16'h241A] = 8'hC5;
DFS[16'h241B] = 8'h4D;
DFS[16'h241C] = 8'h4D;
DFS[16'h241D] = 8'h43;
DFS[16'h241E] = 8'h20;
DFS[16'h241F] = 8'h57;
DFS[16'h2420] = 8'h72;
DFS[16'h2421] = 8'h69;
DFS[16'h2422] = 8'h74;
DFS[16'h2423] = 8'h65;
DFS[16'h2424] = 8'h20;
DFS[16'h2425] = 8'h72;
DFS[16'h2426] = 8'h65;
DFS[16'h2427] = 8'h73;
DFS[16'h2428] = 8'h70;
DFS[16'h2429] = 8'h6F;
DFS[16'h242A] = 8'h6E;
DFS[16'h242B] = 8'h73;
DFS[16'h242C] = 8'h65;
DFS[16'h242D] = 8'h20;
DFS[16'h242E] = 8'h66;
DFS[16'h242F] = 8'h61;
DFS[16'h2430] = 8'h75;
DFS[16'h2431] = 8'h6C;
DFS[16'h2432] = 8'h74;
DFS[16'h2433] = 8'h20;
DFS[16'h2434] = 8'h00;
DFS[16'h2435] = 8'h2C;
DFS[16'h2436] = 8'h40;
DFS[16'h2437] = 8'h0D;
DFS[16'h2438] = 8'h30;
DFS[16'h2439] = 8'h1A;
DFS[16'h243A] = 8'hAC;
DFS[16'h243B] = 8'hD6;
DFS[16'h243C] = 8'h10;
DFS[16'h243D] = 8'hD0;
DFS[16'h243E] = 8'h09;
DFS[16'h243F] = 8'hB1;
DFS[16'h2440] = 8'hA0;
DFS[16'h2441] = 8'h20;
DFS[16'h2442] = 8'hB8;
DFS[16'h2443] = 8'hA1;
DFS[16'h2444] = 8'hC8;
DFS[16'h2445] = 8'hD0;
DFS[16'h2446] = 8'hF8;
DFS[16'h2447] = 8'h60;
DFS[16'h2448] = 8'hA0;
DFS[16'h2449] = 8'h00;
DFS[16'h244A] = 8'hAD;
DFS[16'h244B] = 8'hE5;
DFS[16'h244C] = 8'hFE;
DFS[16'h244D] = 8'h20;
DFS[16'h244E] = 8'hB8;
DFS[16'h244F] = 8'hA1;
DFS[16'h2450] = 8'hC8;
DFS[16'h2451] = 8'hD0;
DFS[16'h2452] = 8'hF7;
DFS[16'h2453] = 8'h60;
DFS[16'h2454] = 8'hAC;
DFS[16'h2455] = 8'hD6;
DFS[16'h2456] = 8'h10;
DFS[16'h2457] = 8'hD0;
DFS[16'h2458] = 8'h09;
DFS[16'h2459] = 8'hB1;
DFS[16'h245A] = 8'hA0;
DFS[16'h245B] = 8'h8D;
DFS[16'h245C] = 8'h18;
DFS[16'h245D] = 8'hFE;
DFS[16'h245E] = 8'hC8;
DFS[16'h245F] = 8'hD0;
DFS[16'h2460] = 8'hF8;
DFS[16'h2461] = 8'h60;
DFS[16'h2462] = 8'hA0;
DFS[16'h2463] = 8'h00;
DFS[16'h2464] = 8'hAD;
DFS[16'h2465] = 8'hE5;
DFS[16'h2466] = 8'hFE;
DFS[16'h2467] = 8'h8D;
DFS[16'h2468] = 8'h18;
DFS[16'h2469] = 8'hFE;
DFS[16'h246A] = 8'h20;
DFS[16'h246B] = 8'h58;
DFS[16'h246C] = 8'hA2;
DFS[16'h246D] = 8'h20;
DFS[16'h246E] = 8'h58;
DFS[16'h246F] = 8'hA2;
DFS[16'h2470] = 8'h20;
DFS[16'h2471] = 8'h58;
DFS[16'h2472] = 8'hA2;
DFS[16'h2473] = 8'hC8;
DFS[16'h2474] = 8'hD0;
DFS[16'h2475] = 8'hEE;
DFS[16'h2476] = 8'h60;
DFS[16'h2477] = 8'h2C;
DFS[16'h2478] = 8'h40;
DFS[16'h2479] = 8'h0D;
DFS[16'h247A] = 8'h30;
DFS[16'h247B] = 8'h0C;
DFS[16'h247C] = 8'hA0;
DFS[16'h247D] = 8'h00;
DFS[16'h247E] = 8'hB9;
DFS[16'h247F] = 8'h00;
DFS[16'h2480] = 8'h0E;
DFS[16'h2481] = 8'h20;
DFS[16'h2482] = 8'hB8;
DFS[16'h2483] = 8'hA1;
DFS[16'h2484] = 8'hC8;
DFS[16'h2485] = 8'hD0;
DFS[16'h2486] = 8'hF7;
DFS[16'h2487] = 8'h60;
DFS[16'h2488] = 8'hA0;
DFS[16'h2489] = 8'h00;
DFS[16'h248A] = 8'hEA;
DFS[16'h248B] = 8'hB9;
DFS[16'h248C] = 8'h00;
DFS[16'h248D] = 8'h0E;
DFS[16'h248E] = 8'h8D;
DFS[16'h248F] = 8'h18;
DFS[16'h2490] = 8'hFE;
DFS[16'h2491] = 8'hC8;
DFS[16'h2492] = 8'hD0;
DFS[16'h2493] = 8'hF6;
DFS[16'h2494] = 8'h60;
DFS[16'h2495] = 8'h9D;
DFS[16'h2496] = 8'h43;
DFS[16'h2497] = 8'h0D;
DFS[16'h2498] = 8'hA9;
DFS[16'h2499] = 8'h00;
DFS[16'h249A] = 8'h9D;
DFS[16'h249B] = 8'h44;
DFS[16'h249C] = 8'h0D;
DFS[16'h249D] = 8'h9D;
DFS[16'h249E] = 8'h45;
DFS[16'h249F] = 8'h0D;
DFS[16'h24A0] = 8'h9D;
DFS[16'h24A1] = 8'h46;
DFS[16'h24A2] = 8'h0D;
DFS[16'h24A3] = 8'h9D;
DFS[16'h24A4] = 8'h47;
DFS[16'h24A5] = 8'h0D;
DFS[16'h24A6] = 8'hA9;
DFS[16'h24A7] = 8'hFF;
DFS[16'h24A8] = 8'h9D;
DFS[16'h24A9] = 8'h42;
DFS[16'h24AA] = 8'h0D;
DFS[16'h24AB] = 8'h9D;
DFS[16'h24AC] = 8'h48;
DFS[16'h24AD] = 8'h0D;
DFS[16'h24AE] = 8'h9D;
DFS[16'h24AF] = 8'h49;
DFS[16'h24B0] = 8'h0D;
DFS[16'h24B1] = 8'hAE;
DFS[16'h24B2] = 8'h03;
DFS[16'h24B3] = 8'h0D;
DFS[16'h24B4] = 8'hBD;
DFS[16'h24B5] = 8'hD2;
DFS[16'h24B6] = 8'hA4;
DFS[16'h24B7] = 8'h8D;
DFS[16'h24B8] = 8'h40;
DFS[16'h24B9] = 8'h0D;
DFS[16'h24BA] = 8'h60;
DFS[16'h24BB] = 8'h2C;
DFS[16'h24BC] = 8'hC9;
DFS[16'h24BD] = 8'h10;
DFS[16'h24BE] = 8'h30;
DFS[16'h24BF] = 8'h11;
DFS[16'h24C0] = 8'hA9;
DFS[16'h24C1] = 8'h8F;
DFS[16'h24C2] = 8'hA2;
DFS[16'h24C3] = 8'h0C;
DFS[16'h24C4] = 8'hA0;
DFS[16'h24C5] = 8'hFF;
DFS[16'h24C6] = 8'h20;
DFS[16'h24C7] = 8'hF4;
DFS[16'h24C8] = 8'hFF;
DFS[16'h24C9] = 8'h8C;
DFS[16'h24CA] = 8'h01;
DFS[16'h24CB] = 8'h0D;
DFS[16'h24CC] = 8'hA9;
DFS[16'h24CD] = 8'hFF;
DFS[16'h24CE] = 8'h8D;
DFS[16'h24CF] = 8'hC9;
DFS[16'h24D0] = 8'h10;
DFS[16'h24D1] = 8'h60;
DFS[16'h24D2] = 8'h80;
DFS[16'h24D3] = 8'h00;
DFS[16'h24D4] = 8'hA9;
DFS[16'h24D5] = 8'h03;
DFS[16'h24D6] = 8'h8D;
DFS[16'h24D7] = 8'h62;
DFS[16'h24D8] = 8'hFE;
DFS[16'h24D9] = 8'hA9;
DFS[16'h24DA] = 8'h00;
DFS[16'h24DB] = 8'h8D;
DFS[16'h24DC] = 8'h60;
DFS[16'h24DD] = 8'hFE;
DFS[16'h24DE] = 8'hAD;
DFS[16'h24DF] = 8'h6B;
DFS[16'h24E0] = 8'hFE;
DFS[16'h24E1] = 8'h29;
DFS[16'h24E2] = 8'hE3;
DFS[16'h24E3] = 8'h8D;
DFS[16'h24E4] = 8'h6B;
DFS[16'h24E5] = 8'hFE;
DFS[16'h24E6] = 8'hA9;
DFS[16'h24E7] = 8'h1C;
DFS[16'h24E8] = 8'h8D;
DFS[16'h24E9] = 8'h6E;
DFS[16'h24EA] = 8'hFE;
DFS[16'h24EB] = 8'h60;
DFS[16'h24EC] = 8'hAD;
DFS[16'h24ED] = 8'h02;
DFS[16'h24EE] = 8'h0D;
DFS[16'h24EF] = 8'hC9;
DFS[16'h24F0] = 8'h54;
DFS[16'h24F1] = 8'hD0;
DFS[16'h24F2] = 8'h04;
DFS[16'h24F3] = 8'h20;
DFS[16'h24F4] = 8'hD4;
DFS[16'h24F5] = 8'hA4;
DFS[16'h24F6] = 8'h60;
DFS[16'h24F7] = 8'h20;
DFS[16'h24F8] = 8'h06;
DFS[16'h24F9] = 8'hA5;
DFS[16'h24FA] = 8'hD0;
DFS[16'h24FB] = 8'hFA;
DFS[16'h24FC] = 8'h20;
DFS[16'h24FD] = 8'h00;
DFS[16'h24FE] = 8'hA0;
DFS[16'h24FF] = 8'hFF;
DFS[16'h2500] = 8'h43;
DFS[16'h2501] = 8'h61;
DFS[16'h2502] = 8'h72;
DFS[16'h2503] = 8'h64;
DFS[16'h2504] = 8'h3F;
DFS[16'h2505] = 8'h00;
DFS[16'h2506] = 8'h20;
DFS[16'h2507] = 8'h71;
DFS[16'h2508] = 8'hA1;
DFS[16'h2509] = 8'hA2;
DFS[16'h250A] = 8'hFF;
DFS[16'h250B] = 8'h8E;
DFS[16'h250C] = 8'h03;
DFS[16'h250D] = 8'h0D;
DFS[16'h250E] = 8'h20;
DFS[16'h250F] = 8'hBB;
DFS[16'h2510] = 8'hA4;
DFS[16'h2511] = 8'hA2;
DFS[16'h2512] = 8'h00;
DFS[16'h2513] = 8'hA9;
DFS[16'h2514] = 8'h40;
DFS[16'h2515] = 8'h20;
DFS[16'h2516] = 8'h95;
DFS[16'h2517] = 8'hA4;
DFS[16'h2518] = 8'hA9;
DFS[16'h2519] = 8'h95;
DFS[16'h251A] = 8'h8D;
DFS[16'h251B] = 8'h48;
DFS[16'h251C] = 8'h0D;
DFS[16'h251D] = 8'hA2;
DFS[16'h251E] = 8'h08;
DFS[16'h251F] = 8'hA9;
DFS[16'h2520] = 8'h41;
DFS[16'h2521] = 8'h20;
DFS[16'h2522] = 8'h95;
DFS[16'h2523] = 8'hA4;
DFS[16'h2524] = 8'h20;
DFS[16'h2525] = 8'hD4;
DFS[16'h2526] = 8'hA4;
DFS[16'h2527] = 8'hA9;
DFS[16'h2528] = 8'h32;
DFS[16'h2529] = 8'h85;
DFS[16'h252A] = 8'hA6;
DFS[16'h252B] = 8'hAE;
DFS[16'h252C] = 8'h04;
DFS[16'h252D] = 8'h0D;
DFS[16'h252E] = 8'hE0;
DFS[16'h252F] = 8'h02;
DFS[16'h2530] = 8'hB0;
DFS[16'h2531] = 8'h5A;
DFS[16'h2532] = 8'h8E;
DFS[16'h2533] = 8'h03;
DFS[16'h2534] = 8'h0D;
DFS[16'h2535] = 8'hBD;
DFS[16'h2536] = 8'hD2;
DFS[16'h2537] = 8'hA4;
DFS[16'h2538] = 8'h8D;
DFS[16'h2539] = 8'h40;
DFS[16'h253A] = 8'h0D;
DFS[16'h253B] = 8'hA0;
DFS[16'h253C] = 8'h0A;
DFS[16'h253D] = 8'h20;
DFS[16'h253E] = 8'h10;
DFS[16'h253F] = 8'hA2;
DFS[16'h2540] = 8'hA2;
DFS[16'h2541] = 8'h00;
DFS[16'h2542] = 8'h20;
DFS[16'h2543] = 8'h59;
DFS[16'h2544] = 8'hA2;
DFS[16'h2545] = 8'h29;
DFS[16'h2546] = 8'h81;
DFS[16'h2547] = 8'hC9;
DFS[16'h2548] = 8'h01;
DFS[16'h2549] = 8'hD0;
DFS[16'h254A] = 8'h35;
DFS[16'h254B] = 8'h24;
DFS[16'h254C] = 8'hFF;
DFS[16'h254D] = 8'h30;
DFS[16'h254E] = 8'h31;
DFS[16'h254F] = 8'hA2;
DFS[16'h2550] = 8'h08;
DFS[16'h2551] = 8'h20;
DFS[16'h2552] = 8'h59;
DFS[16'h2553] = 8'hA2;
DFS[16'h2554] = 8'hC9;
DFS[16'h2555] = 8'h02;
DFS[16'h2556] = 8'hB0;
DFS[16'h2557] = 8'h28;
DFS[16'h2558] = 8'hC9;
DFS[16'h2559] = 8'h00;
DFS[16'h255A] = 8'hD0;
DFS[16'h255B] = 8'hEF;
DFS[16'h255C] = 8'hA2;
DFS[16'h255D] = 8'h00;
DFS[16'h255E] = 8'hA9;
DFS[16'h255F] = 8'h50;
DFS[16'h2560] = 8'h20;
DFS[16'h2561] = 8'h95;
DFS[16'h2562] = 8'hA4;
DFS[16'h2563] = 8'hA9;
DFS[16'h2564] = 8'h02;
DFS[16'h2565] = 8'h8D;
DFS[16'h2566] = 8'h46;
DFS[16'h2567] = 8'h0D;
DFS[16'h2568] = 8'hA2;
DFS[16'h2569] = 8'h00;
DFS[16'h256A] = 8'h20;
DFS[16'h256B] = 8'h59;
DFS[16'h256C] = 8'hA2;
DFS[16'h256D] = 8'hD0;
DFS[16'h256E] = 8'h23;
DFS[16'h256F] = 8'hA9;
DFS[16'h2570] = 8'h54;
DFS[16'h2571] = 8'h8D;
DFS[16'h2572] = 8'h02;
DFS[16'h2573] = 8'h0D;
DFS[16'h2574] = 8'hAD;
DFS[16'h2575] = 8'h03;
DFS[16'h2576] = 8'h0D;
DFS[16'h2577] = 8'h8D;
DFS[16'h2578] = 8'h04;
DFS[16'h2579] = 8'h0D;
DFS[16'h257A] = 8'h20;
DFS[16'h257B] = 8'h7B;
DFS[16'h257C] = 8'hA1;
DFS[16'h257D] = 8'hA9;
DFS[16'h257E] = 8'hFF;
DFS[16'h257F] = 8'h60;
DFS[16'h2580] = 8'hAE;
DFS[16'h2581] = 8'h03;
DFS[16'h2582] = 8'h0D;
DFS[16'h2583] = 8'hE8;
DFS[16'h2584] = 8'hE0;
DFS[16'h2585] = 8'h02;
DFS[16'h2586] = 8'h90;
DFS[16'h2587] = 8'hAA;
DFS[16'h2588] = 8'hC6;
DFS[16'h2589] = 8'hA6;
DFS[16'h258A] = 8'hD0;
DFS[16'h258B] = 8'h9F;
DFS[16'h258C] = 8'hA9;
DFS[16'h258D] = 8'h00;
DFS[16'h258E] = 8'h8D;
DFS[16'h258F] = 8'h02;
DFS[16'h2590] = 8'h0D;
DFS[16'h2591] = 8'h60;
DFS[16'h2592] = 8'h20;
DFS[16'h2593] = 8'h1F;
DFS[16'h2594] = 8'hA0;
DFS[16'h2595] = 8'hFF;
DFS[16'h2596] = 8'h53;
DFS[16'h2597] = 8'h65;
DFS[16'h2598] = 8'h74;
DFS[16'h2599] = 8'h20;
DFS[16'h259A] = 8'h62;
DFS[16'h259B] = 8'h6C;
DFS[16'h259C] = 8'h6F;
DFS[16'h259D] = 8'h63;
DFS[16'h259E] = 8'h6B;
DFS[16'h259F] = 8'h20;
DFS[16'h25A0] = 8'h6C;
DFS[16'h25A1] = 8'h65;
DFS[16'h25A2] = 8'h6E;
DFS[16'h25A3] = 8'h20;
DFS[16'h25A4] = 8'h65;
DFS[16'h25A5] = 8'h72;
DFS[16'h25A6] = 8'h72;
DFS[16'h25A7] = 8'h6F;
DFS[16'h25A8] = 8'h72;
DFS[16'h25A9] = 8'h20;
DFS[16'h25AA] = 8'h00;
DFS[16'h25AB] = 8'hA9;
DFS[16'h25AC] = 8'h51;
DFS[16'h25AD] = 8'hA2;
DFS[16'h25AE] = 8'h00;
DFS[16'h25AF] = 8'h20;
DFS[16'h25B0] = 8'h95;
DFS[16'h25B1] = 8'hA4;
DFS[16'h25B2] = 8'hA5;
DFS[16'h25B3] = 8'hA2;
DFS[16'h25B4] = 8'h8D;
DFS[16'h25B5] = 8'h46;
DFS[16'h25B6] = 8'h0D;
DFS[16'h25B7] = 8'hA5;
DFS[16'h25B8] = 8'hA3;
DFS[16'h25B9] = 8'h8D;
DFS[16'h25BA] = 8'h45;
DFS[16'h25BB] = 8'h0D;
DFS[16'h25BC] = 8'hA5;
DFS[16'h25BD] = 8'hA4;
DFS[16'h25BE] = 8'h8D;
DFS[16'h25BF] = 8'h44;
DFS[16'h25C0] = 8'h0D;
DFS[16'h25C1] = 8'h60;
DFS[16'h25C2] = 8'hA2;
DFS[16'h25C3] = 8'h00;
DFS[16'h25C4] = 8'h20;
DFS[16'h25C5] = 8'h59;
DFS[16'h25C6] = 8'hA2;
DFS[16'h25C7] = 8'hD0;
DFS[16'h25C8] = 8'h04;
DFS[16'h25C9] = 8'h20;
DFS[16'h25CA] = 8'hB6;
DFS[16'h25CB] = 8'hA2;
DFS[16'h25CC] = 8'h60;
DFS[16'h25CD] = 8'h20;
DFS[16'h25CE] = 8'h1F;
DFS[16'h25CF] = 8'hA0;
DFS[16'h25D0] = 8'hC5;
DFS[16'h25D1] = 8'h4D;
DFS[16'h25D2] = 8'h4D;
DFS[16'h25D3] = 8'h43;
DFS[16'h25D4] = 8'h20;
DFS[16'h25D5] = 8'h52;
DFS[16'h25D6] = 8'h65;
DFS[16'h25D7] = 8'h61;
DFS[16'h25D8] = 8'h64;
DFS[16'h25D9] = 8'h20;
DFS[16'h25DA] = 8'h66;
DFS[16'h25DB] = 8'h61;
DFS[16'h25DC] = 8'h75;
DFS[16'h25DD] = 8'h6C;
DFS[16'h25DE] = 8'h74;
DFS[16'h25DF] = 8'h20;
DFS[16'h25E0] = 8'h00;
DFS[16'h25E1] = 8'hA2;
DFS[16'h25E2] = 8'h00;
DFS[16'h25E3] = 8'h20;
DFS[16'h25E4] = 8'h59;
DFS[16'h25E5] = 8'hA2;
DFS[16'h25E6] = 8'hD0;
DFS[16'h25E7] = 8'h03;
DFS[16'h25E8] = 8'h4C;
DFS[16'h25E9] = 8'hB0;
DFS[16'h25EA] = 8'hA3;
DFS[16'h25EB] = 8'h20;
DFS[16'h25EC] = 8'h1F;
DFS[16'h25ED] = 8'hA0;
DFS[16'h25EE] = 8'hC5;
DFS[16'h25EF] = 8'h4D;
DFS[16'h25F0] = 8'h4D;
DFS[16'h25F1] = 8'h43;
DFS[16'h25F2] = 8'h20;
DFS[16'h25F3] = 8'h57;
DFS[16'h25F4] = 8'h72;
DFS[16'h25F5] = 8'h69;
DFS[16'h25F6] = 8'h74;
DFS[16'h25F7] = 8'h65;
DFS[16'h25F8] = 8'h20;
DFS[16'h25F9] = 8'h66;
DFS[16'h25FA] = 8'h61;
DFS[16'h25FB] = 8'h75;
DFS[16'h25FC] = 8'h6C;
DFS[16'h25FD] = 8'h74;
DFS[16'h25FE] = 8'h20;
DFS[16'h25FF] = 8'h00;
DFS[16'h2600] = 8'h20;
DFS[16'h2601] = 8'h71;
DFS[16'h2602] = 8'hA1;
DFS[16'h2603] = 8'hA9;
DFS[16'h2604] = 8'h00;
DFS[16'h2605] = 8'h8D;
DFS[16'h2606] = 8'hD6;
DFS[16'h2607] = 8'h10;
DFS[16'h2608] = 8'h85;
DFS[16'h2609] = 8'hA0;
DFS[16'h260A] = 8'hA9;
DFS[16'h260B] = 8'h0E;
DFS[16'h260C] = 8'h85;
DFS[16'h260D] = 8'hA1;
DFS[16'h260E] = 8'h60;
DFS[16'h260F] = 8'h20;
DFS[16'h2610] = 8'h00;
DFS[16'h2611] = 8'hA6;
DFS[16'h2612] = 8'h20;
DFS[16'h2613] = 8'hAB;
DFS[16'h2614] = 8'hA5;
DFS[16'h2615] = 8'h20;
DFS[16'h2616] = 8'hC2;
DFS[16'h2617] = 8'hA5;
DFS[16'h2618] = 8'h20;
DFS[16'h2619] = 8'hD5;
DFS[16'h261A] = 8'hA2;
DFS[16'h261B] = 8'hE6;
DFS[16'h261C] = 8'hA1;
DFS[16'h261D] = 8'h20;
DFS[16'h261E] = 8'hD5;
DFS[16'h261F] = 8'hA2;
DFS[16'h2620] = 8'hA0;
DFS[16'h2621] = 8'h02;
DFS[16'h2622] = 8'h20;
DFS[16'h2623] = 8'h10;
DFS[16'h2624] = 8'hA2;
DFS[16'h2625] = 8'h4C;
DFS[16'h2626] = 8'h7B;
DFS[16'h2627] = 8'hA1;
DFS[16'h2628] = 8'h20;
DFS[16'h2629] = 8'h00;
DFS[16'h262A] = 8'hA6;
DFS[16'h262B] = 8'hA9;
DFS[16'h262C] = 8'h58;
DFS[16'h262D] = 8'h20;
DFS[16'h262E] = 8'hAD;
DFS[16'h262F] = 8'hA5;
DFS[16'h2630] = 8'h20;
DFS[16'h2631] = 8'hE1;
DFS[16'h2632] = 8'hA5;
DFS[16'h2633] = 8'h20;
DFS[16'h2634] = 8'h35;
DFS[16'h2635] = 8'hA4;
DFS[16'h2636] = 8'hE6;
DFS[16'h2637] = 8'hA1;
DFS[16'h2638] = 8'h20;
DFS[16'h2639] = 8'h35;
DFS[16'h263A] = 8'hA4;
DFS[16'h263B] = 8'h20;
DFS[16'h263C] = 8'hD2;
DFS[16'h263D] = 8'hA3;
DFS[16'h263E] = 8'h4C;
DFS[16'h263F] = 8'h7B;
DFS[16'h2640] = 8'hA1;
DFS[16'h2641] = 8'h60;
DFS[16'h2642] = 8'h20;
DFS[16'h2643] = 8'h71;
DFS[16'h2644] = 8'hA1;
DFS[16'h2645] = 8'h20;
DFS[16'h2646] = 8'h4B;
DFS[16'h2647] = 8'hA6;
DFS[16'h2648] = 8'h4C;
DFS[16'h2649] = 8'h7B;
DFS[16'h264A] = 8'hA1;
DFS[16'h264B] = 8'hA6;
DFS[16'h264C] = 8'hA5;
DFS[16'h264D] = 8'hF0;
DFS[16'h264E] = 8'hF2;
DFS[16'h264F] = 8'hA9;
DFS[16'h2650] = 8'h01;
DFS[16'h2651] = 8'h20;
DFS[16'h2652] = 8'h98;
DFS[16'h2653] = 8'hA0;
DFS[16'h2654] = 8'hA6;
DFS[16'h2655] = 8'hA5;
DFS[16'h2656] = 8'h66;
DFS[16'h2657] = 8'hA2;
DFS[16'h2658] = 8'h66;
DFS[16'h2659] = 8'hA6;
DFS[16'h265A] = 8'h10;
DFS[16'h265B] = 8'h01;
DFS[16'h265C] = 8'hE8;
DFS[16'h265D] = 8'h86;
DFS[16'h265E] = 8'hA5;
DFS[16'h265F] = 8'h06;
DFS[16'h2660] = 8'hA2;
DFS[16'h2661] = 8'h20;
DFS[16'h2662] = 8'hAB;
DFS[16'h2663] = 8'hA5;
DFS[16'h2664] = 8'hA6;
DFS[16'h2665] = 8'hA5;
DFS[16'h2666] = 8'hE0;
DFS[16'h2667] = 8'h03;
DFS[16'h2668] = 8'hB0;
DFS[16'h2669] = 8'h08;
DFS[16'h266A] = 8'hA5;
DFS[16'h266B] = 8'hA7;
DFS[16'h266C] = 8'hD0;
DFS[16'h266D] = 8'h4F;
DFS[16'h266E] = 8'hE0;
DFS[16'h266F] = 8'h01;
DFS[16'h2670] = 8'hF0;
DFS[16'h2671] = 8'h42;
DFS[16'h2672] = 8'h24;
DFS[16'h2673] = 8'hA6;
DFS[16'h2674] = 8'h10;
DFS[16'h2675] = 8'h0D;
DFS[16'h2676] = 8'h20;
DFS[16'h2677] = 8'hC2;
DFS[16'h2678] = 8'hA5;
DFS[16'h2679] = 8'hA0;
DFS[16'h267A] = 8'h00;
DFS[16'h267B] = 8'h84;
DFS[16'h267C] = 8'hA6;
DFS[16'h267D] = 8'h20;
DFS[16'h267E] = 8'h10;
DFS[16'h267F] = 8'hA2;
DFS[16'h2680] = 8'h4C;
DFS[16'h2681] = 8'h8B;
DFS[16'h2682] = 8'hA6;
DFS[16'h2683] = 8'h20;
DFS[16'h2684] = 8'hC2;
DFS[16'h2685] = 8'hA5;
DFS[16'h2686] = 8'h20;
DFS[16'h2687] = 8'hD5;
DFS[16'h2688] = 8'hA2;
DFS[16'h2689] = 8'hE6;
DFS[16'h268A] = 8'hA1;
DFS[16'h268B] = 8'h20;
DFS[16'h268C] = 8'hD5;
DFS[16'h268D] = 8'hA2;
DFS[16'h268E] = 8'hE6;
DFS[16'h268F] = 8'hA1;
DFS[16'h2690] = 8'hA0;
DFS[16'h2691] = 8'h02;
DFS[16'h2692] = 8'h20;
DFS[16'h2693] = 8'h10;
DFS[16'h2694] = 8'hA2;
DFS[16'h2695] = 8'hEE;
DFS[16'h2696] = 8'h46;
DFS[16'h2697] = 8'h0D;
DFS[16'h2698] = 8'hEE;
DFS[16'h2699] = 8'h46;
DFS[16'h269A] = 8'h0D;
DFS[16'h269B] = 8'hD0;
DFS[16'h269C] = 8'h08;
DFS[16'h269D] = 8'hEE;
DFS[16'h269E] = 8'h45;
DFS[16'h269F] = 8'h0D;
DFS[16'h26A0] = 8'hD0;
DFS[16'h26A1] = 8'h03;
DFS[16'h26A2] = 8'hEE;
DFS[16'h26A3] = 8'h44;
DFS[16'h26A4] = 8'h0D;
DFS[16'h26A5] = 8'hA6;
DFS[16'h26A6] = 8'hA5;
DFS[16'h26A7] = 8'hCA;
DFS[16'h26A8] = 8'hCA;
DFS[16'h26A9] = 8'hF0;
DFS[16'h26AA] = 8'h96;
DFS[16'h26AB] = 8'h86;
DFS[16'h26AC] = 8'hA5;
DFS[16'h26AD] = 8'hE0;
DFS[16'h26AE] = 8'h03;
DFS[16'h26AF] = 8'hB0;
DFS[16'h26B0] = 8'hD2;
DFS[16'h26B1] = 8'h4C;
DFS[16'h26B2] = 8'h6A;
DFS[16'h26B3] = 8'hA6;
DFS[16'h26B4] = 8'h20;
DFS[16'h26B5] = 8'hC2;
DFS[16'h26B6] = 8'hA5;
DFS[16'h26B7] = 8'h20;
DFS[16'h26B8] = 8'hD5;
DFS[16'h26B9] = 8'hA2;
DFS[16'h26BA] = 8'h4C;
DFS[16'h26BB] = 8'hE4;
DFS[16'h26BC] = 8'hA6;
DFS[16'h26BD] = 8'h20;
DFS[16'h26BE] = 8'hC2;
DFS[16'h26BF] = 8'hA5;
DFS[16'h26C0] = 8'h24;
DFS[16'h26C1] = 8'hA6;
DFS[16'h26C2] = 8'h10;
DFS[16'h26C3] = 8'h08;
DFS[16'h26C4] = 8'hA0;
DFS[16'h26C5] = 8'h00;
DFS[16'h26C6] = 8'h20;
DFS[16'h26C7] = 8'h10;
DFS[16'h26C8] = 8'hA2;
DFS[16'h26C9] = 8'h4C;
DFS[16'h26CA] = 8'hD5;
DFS[16'h26CB] = 8'hA6;
DFS[16'h26CC] = 8'hC6;
DFS[16'h26CD] = 8'hA5;
DFS[16'h26CE] = 8'hF0;
DFS[16'h26CF] = 8'h05;
DFS[16'h26D0] = 8'h20;
DFS[16'h26D1] = 8'hD5;
DFS[16'h26D2] = 8'hA2;
DFS[16'h26D3] = 8'hE6;
DFS[16'h26D4] = 8'hA1;
DFS[16'h26D5] = 8'h20;
DFS[16'h26D6] = 8'h14;
DFS[16'h26D7] = 8'hA3;
DFS[16'h26D8] = 8'h98;
DFS[16'h26D9] = 8'h49;
DFS[16'h26DA] = 8'hFF;
DFS[16'h26DB] = 8'hA8;
DFS[16'h26DC] = 8'hC8;
DFS[16'h26DD] = 8'h20;
DFS[16'h26DE] = 8'h10;
DFS[16'h26DF] = 8'hA2;
DFS[16'h26E0] = 8'hA5;
DFS[16'h26E1] = 8'hA5;
DFS[16'h26E2] = 8'hD0;
DFS[16'h26E3] = 8'h05;
DFS[16'h26E4] = 8'hA0;
DFS[16'h26E5] = 8'h00;
DFS[16'h26E6] = 8'h20;
DFS[16'h26E7] = 8'h10;
DFS[16'h26E8] = 8'hA2;
DFS[16'h26E9] = 8'hA0;
DFS[16'h26EA] = 8'h02;
DFS[16'h26EB] = 8'h4C;
DFS[16'h26EC] = 8'h10;
DFS[16'h26ED] = 8'hA2;
DFS[16'h26EE] = 8'h60;
DFS[16'h26EF] = 8'h20;
DFS[16'h26F0] = 8'h71;
DFS[16'h26F1] = 8'hA1;
DFS[16'h26F2] = 8'h20;
DFS[16'h26F3] = 8'hF8;
DFS[16'h26F4] = 8'hA6;
DFS[16'h26F5] = 8'h4C;
DFS[16'h26F6] = 8'h7B;
DFS[16'h26F7] = 8'hA1;
DFS[16'h26F8] = 8'hA6;
DFS[16'h26F9] = 8'hA5;
DFS[16'h26FA] = 8'hF0;
DFS[16'h26FB] = 8'hF2;
DFS[16'h26FC] = 8'hA9;
DFS[16'h26FD] = 8'h00;
DFS[16'h26FE] = 8'h20;
DFS[16'h26FF] = 8'h98;
DFS[16'h2700] = 8'hA0;
DFS[16'h2701] = 8'hA6;
DFS[16'h2702] = 8'hA5;
DFS[16'h2703] = 8'h66;
DFS[16'h2704] = 8'hA2;
DFS[16'h2705] = 8'h6A;
DFS[16'h2706] = 8'h06;
DFS[16'h2707] = 8'hA2;
DFS[16'h2708] = 8'h48;
DFS[16'h2709] = 8'hA9;
DFS[16'h270A] = 8'h58;
DFS[16'h270B] = 8'h20;
DFS[16'h270C] = 8'hAD;
DFS[16'h270D] = 8'hA5;
DFS[16'h270E] = 8'h68;
DFS[16'h270F] = 8'h10;
DFS[16'h2710] = 8'h41;
DFS[16'h2711] = 8'hA9;
DFS[16'h2712] = 8'hFF;
DFS[16'h2713] = 8'h8D;
DFS[16'h2714] = 8'h82;
DFS[16'h2715] = 8'h10;
DFS[16'h2716] = 8'hA9;
DFS[16'h2717] = 8'h51;
DFS[16'h2718] = 8'h8D;
DFS[16'h2719] = 8'h43;
DFS[16'h271A] = 8'h0D;
DFS[16'h271B] = 8'h20;
DFS[16'h271C] = 8'hC2;
DFS[16'h271D] = 8'hA5;
DFS[16'h271E] = 8'h20;
DFS[16'h271F] = 8'h7E;
DFS[16'h2720] = 8'hA3;
DFS[16'h2721] = 8'hA0;
DFS[16'h2722] = 8'h00;
DFS[16'h2723] = 8'h20;
DFS[16'h2724] = 8'h10;
DFS[16'h2725] = 8'hA2;
DFS[16'h2726] = 8'hA0;
DFS[16'h2727] = 8'h02;
DFS[16'h2728] = 8'h20;
DFS[16'h2729] = 8'h10;
DFS[16'h272A] = 8'hA2;
DFS[16'h272B] = 8'hA9;
DFS[16'h272C] = 8'h58;
DFS[16'h272D] = 8'h8D;
DFS[16'h272E] = 8'h43;
DFS[16'h272F] = 8'h0D;
DFS[16'h2730] = 8'h20;
DFS[16'h2731] = 8'hE1;
DFS[16'h2732] = 8'hA5;
DFS[16'h2733] = 8'h20;
DFS[16'h2734] = 8'h77;
DFS[16'h2735] = 8'hA4;
DFS[16'h2736] = 8'h20;
DFS[16'h2737] = 8'h35;
DFS[16'h2738] = 8'hA4;
DFS[16'h2739] = 8'h20;
DFS[16'h273A] = 8'hD2;
DFS[16'h273B] = 8'hA3;
DFS[16'h273C] = 8'hC6;
DFS[16'h273D] = 8'hA5;
DFS[16'h273E] = 8'hF0;
DFS[16'h273F] = 8'hAE;
DFS[16'h2740] = 8'hE6;
DFS[16'h2741] = 8'hA1;
DFS[16'h2742] = 8'hEE;
DFS[16'h2743] = 8'h46;
DFS[16'h2744] = 8'h0D;
DFS[16'h2745] = 8'hEE;
DFS[16'h2746] = 8'h46;
DFS[16'h2747] = 8'h0D;
DFS[16'h2748] = 8'hD0;
DFS[16'h2749] = 8'h08;
DFS[16'h274A] = 8'hEE;
DFS[16'h274B] = 8'h45;
DFS[16'h274C] = 8'h0D;
DFS[16'h274D] = 8'hD0;
DFS[16'h274E] = 8'h03;
DFS[16'h274F] = 8'hEE;
DFS[16'h2750] = 8'h44;
DFS[16'h2751] = 8'h0D;
DFS[16'h2752] = 8'hA6;
DFS[16'h2753] = 8'hA5;
DFS[16'h2754] = 8'hF0;
DFS[16'h2755] = 8'h44;
DFS[16'h2756] = 8'hCA;
DFS[16'h2757] = 8'hD0;
DFS[16'h2758] = 8'h2B;
DFS[16'h2759] = 8'hA9;
DFS[16'h275A] = 8'hFF;
DFS[16'h275B] = 8'h8D;
DFS[16'h275C] = 8'h82;
DFS[16'h275D] = 8'h10;
DFS[16'h275E] = 8'hA9;
DFS[16'h275F] = 8'h51;
DFS[16'h2760] = 8'h8D;
DFS[16'h2761] = 8'h43;
DFS[16'h2762] = 8'h0D;
DFS[16'h2763] = 8'h20;
DFS[16'h2764] = 8'hC2;
DFS[16'h2765] = 8'hA5;
DFS[16'h2766] = 8'hA0;
DFS[16'h2767] = 8'h00;
DFS[16'h2768] = 8'h20;
DFS[16'h2769] = 8'h10;
DFS[16'h276A] = 8'hA2;
DFS[16'h276B] = 8'h20;
DFS[16'h276C] = 8'h7E;
DFS[16'h276D] = 8'hA3;
DFS[16'h276E] = 8'hA0;
DFS[16'h276F] = 8'h02;
DFS[16'h2770] = 8'h20;
DFS[16'h2771] = 8'h10;
DFS[16'h2772] = 8'hA2;
DFS[16'h2773] = 8'hA9;
DFS[16'h2774] = 8'h58;
DFS[16'h2775] = 8'h8D;
DFS[16'h2776] = 8'h43;
DFS[16'h2777] = 8'h0D;
DFS[16'h2778] = 8'h20;
DFS[16'h2779] = 8'hE1;
DFS[16'h277A] = 8'hA5;
DFS[16'h277B] = 8'h20;
DFS[16'h277C] = 8'h35;
DFS[16'h277D] = 8'hA4;
DFS[16'h277E] = 8'h20;
DFS[16'h277F] = 8'h77;
DFS[16'h2780] = 8'hA4;
DFS[16'h2781] = 8'h4C;
DFS[16'h2782] = 8'hD2;
DFS[16'h2783] = 8'hA3;
DFS[16'h2784] = 8'h20;
DFS[16'h2785] = 8'hE1;
DFS[16'h2786] = 8'hA5;
DFS[16'h2787] = 8'h20;
DFS[16'h2788] = 8'h35;
DFS[16'h2789] = 8'hA4;
DFS[16'h278A] = 8'hE6;
DFS[16'h278B] = 8'hA1;
DFS[16'h278C] = 8'h20;
DFS[16'h278D] = 8'h35;
DFS[16'h278E] = 8'hA4;
DFS[16'h278F] = 8'hE6;
DFS[16'h2790] = 8'hA1;
DFS[16'h2791] = 8'h20;
DFS[16'h2792] = 8'hD2;
DFS[16'h2793] = 8'hA3;
DFS[16'h2794] = 8'hC6;
DFS[16'h2795] = 8'hA5;
DFS[16'h2796] = 8'hC6;
DFS[16'h2797] = 8'hA5;
DFS[16'h2798] = 8'hD0;
DFS[16'h2799] = 8'hA8;
DFS[16'h279A] = 8'h60;
DFS[16'h279B] = 8'hA9;
DFS[16'h279C] = 8'h51;
DFS[16'h279D] = 8'hA2;
DFS[16'h279E] = 8'h08;
DFS[16'h279F] = 8'h20;
DFS[16'h27A0] = 8'h95;
DFS[16'h27A1] = 8'hA4;
DFS[16'h27A2] = 8'hA5;
DFS[16'h27A3] = 8'hA2;
DFS[16'h27A4] = 8'h8D;
DFS[16'h27A5] = 8'h4E;
DFS[16'h27A6] = 8'h0D;
DFS[16'h27A7] = 8'hA5;
DFS[16'h27A8] = 8'hA3;
DFS[16'h27A9] = 8'h8D;
DFS[16'h27AA] = 8'h4D;
DFS[16'h27AB] = 8'h0D;
DFS[16'h27AC] = 8'hA5;
DFS[16'h27AD] = 8'hA4;
DFS[16'h27AE] = 8'h8D;
DFS[16'h27AF] = 8'h4C;
DFS[16'h27B0] = 8'h0D;
DFS[16'h27B1] = 8'h60;
DFS[16'h27B2] = 8'h20;
DFS[16'h27B3] = 8'h71;
DFS[16'h27B4] = 8'hA1;
DFS[16'h27B5] = 8'hA2;
DFS[16'h27B6] = 8'h08;
DFS[16'h27B7] = 8'h20;
DFS[16'h27B8] = 8'hC4;
DFS[16'h27B9] = 8'hA5;
DFS[16'h27BA] = 8'hA9;
DFS[16'h27BB] = 8'h5F;
DFS[16'h27BC] = 8'h85;
DFS[16'h27BD] = 8'hA0;
DFS[16'h27BE] = 8'hA9;
DFS[16'h27BF] = 8'h0D;
DFS[16'h27C0] = 8'h85;
DFS[16'h27C1] = 8'hA1;
DFS[16'h27C2] = 8'hA9;
DFS[16'h27C3] = 8'h08;
DFS[16'h27C4] = 8'h85;
DFS[16'h27C5] = 8'hA7;
DFS[16'h27C6] = 8'h20;
DFS[16'h27C7] = 8'h14;
DFS[16'h27C8] = 8'hA3;
DFS[16'h27C9] = 8'hA0;
DFS[16'h27CA] = 8'hF8;
DFS[16'h27CB] = 8'h20;
DFS[16'h27CC] = 8'h10;
DFS[16'h27CD] = 8'hA2;
DFS[16'h27CE] = 8'hA9;
DFS[16'h27CF] = 8'h67;
DFS[16'h27D0] = 8'h85;
DFS[16'h27D1] = 8'hA0;
DFS[16'h27D2] = 8'hA9;
DFS[16'h27D3] = 8'h08;
DFS[16'h27D4] = 8'h85;
DFS[16'h27D5] = 8'hA7;
DFS[16'h27D6] = 8'h20;
DFS[16'h27D7] = 8'h14;
DFS[16'h27D8] = 8'hA3;
DFS[16'h27D9] = 8'hA0;
DFS[16'h27DA] = 8'hFA;
DFS[16'h27DB] = 8'h20;
DFS[16'h27DC] = 8'h10;
DFS[16'h27DD] = 8'hA2;
DFS[16'h27DE] = 8'h18;
DFS[16'h27DF] = 8'hAD;
DFS[16'h27E0] = 8'h4E;
DFS[16'h27E1] = 8'h0D;
DFS[16'h27E2] = 8'h69;
DFS[16'h27E3] = 8'h20;
DFS[16'h27E4] = 8'h8D;
DFS[16'h27E5] = 8'h4E;
DFS[16'h27E6] = 8'h0D;
DFS[16'h27E7] = 8'hAD;
DFS[16'h27E8] = 8'h4D;
DFS[16'h27E9] = 8'h0D;
DFS[16'h27EA] = 8'h69;
DFS[16'h27EB] = 8'h03;
DFS[16'h27EC] = 8'h8D;
DFS[16'h27ED] = 8'h4D;
DFS[16'h27EE] = 8'h0D;
DFS[16'h27EF] = 8'h90;
DFS[16'h27F0] = 8'h03;
DFS[16'h27F1] = 8'hEE;
DFS[16'h27F2] = 8'h4C;
DFS[16'h27F3] = 8'h0D;
DFS[16'h27F4] = 8'h4C;
DFS[16'h27F5] = 8'h7B;
DFS[16'h27F6] = 8'hA1;
DFS[16'h27F7] = 8'h20;
DFS[16'h27F8] = 8'h06;
DFS[16'h27F9] = 8'hA5;
DFS[16'h27FA] = 8'hF0;
DFS[16'h27FB] = 8'hB5;
DFS[16'h27FC] = 8'hA9;
DFS[16'h27FD] = 8'h7A;
DFS[16'h27FE] = 8'h20;
DFS[16'h27FF] = 8'hF4;
DFS[16'h2800] = 8'hFF;
DFS[16'h2801] = 8'h8A;
DFS[16'h2802] = 8'h30;
DFS[16'h2803] = 8'h0D;
DFS[16'h2804] = 8'hC9;
DFS[16'h2805] = 8'h65;
DFS[16'h2806] = 8'hF0;
DFS[16'h2807] = 8'h04;
DFS[16'h2808] = 8'hC9;
DFS[16'h2809] = 8'h42;
DFS[16'h280A] = 8'hD0;
DFS[16'h280B] = 8'hA5;
DFS[16'h280C] = 8'hA9;
DFS[16'h280D] = 8'h78;
DFS[16'h280E] = 8'h20;
DFS[16'h280F] = 8'hF4;
DFS[16'h2810] = 8'hFF;
DFS[16'h2811] = 8'h8E;
DFS[16'h2812] = 8'h52;
DFS[16'h2813] = 8'h0D;
DFS[16'h2814] = 8'h4C;
DFS[16'h2815] = 8'h20;
DFS[16'h2816] = 8'h93;
DFS[16'h2817] = 8'hAD;
DFS[16'h2818] = 8'h05;
DFS[16'h2819] = 8'h0D;
DFS[16'h281A] = 8'hC9;
DFS[16'h281B] = 8'h54;
DFS[16'h281C] = 8'hD0;
DFS[16'h281D] = 8'h17;
DFS[16'h281E] = 8'hAD;
DFS[16'h281F] = 8'h06;
DFS[16'h2820] = 8'h0D;
DFS[16'h2821] = 8'h4D;
DFS[16'h2822] = 8'h09;
DFS[16'h2823] = 8'h0D;
DFS[16'h2824] = 8'h4D;
DFS[16'h2825] = 8'h07;
DFS[16'h2826] = 8'h0D;
DFS[16'h2827] = 8'h4D;
DFS[16'h2828] = 8'h0A;
DFS[16'h2829] = 8'h0D;
DFS[16'h282A] = 8'h4D;
DFS[16'h282B] = 8'h08;
DFS[16'h282C] = 8'h0D;
DFS[16'h282D] = 8'h4D;
DFS[16'h282E] = 8'h0B;
DFS[16'h282F] = 8'h0D;
DFS[16'h2830] = 8'hC9;
DFS[16'h2831] = 8'hFF;
DFS[16'h2832] = 8'hD0;
DFS[16'h2833] = 8'h01;
DFS[16'h2834] = 8'h60;
DFS[16'h2835] = 8'hA2;
DFS[16'h2836] = 8'h08;
DFS[16'h2837] = 8'hB5;
DFS[16'h2838] = 8'hA1;
DFS[16'h2839] = 8'h48;
DFS[16'h283A] = 8'hCA;
DFS[16'h283B] = 8'hD0;
DFS[16'h283C] = 8'hFA;
DFS[16'h283D] = 8'hA9;
DFS[16'h283E] = 8'h00;
DFS[16'h283F] = 8'h85;
DFS[16'h2840] = 8'hA2;
DFS[16'h2841] = 8'h85;
DFS[16'h2842] = 8'hA3;
DFS[16'h2843] = 8'h85;
DFS[16'h2844] = 8'hA4;
DFS[16'h2845] = 8'h20;
DFS[16'h2846] = 8'h0F;
DFS[16'h2847] = 8'hA6;
DFS[16'h2848] = 8'hA9;
DFS[16'h2849] = 8'hDD;
DFS[16'h284A] = 8'h8D;
DFS[16'h284B] = 8'h82;
DFS[16'h284C] = 8'h10;
DFS[16'h284D] = 8'h20;
DFS[16'h284E] = 8'h6B;
DFS[16'h284F] = 8'hA8;
DFS[16'h2850] = 8'hF0;
DFS[16'h2851] = 8'h29;
DFS[16'h2852] = 8'hA9;
DFS[16'h2853] = 8'h00;
DFS[16'h2854] = 8'h8D;
DFS[16'h2855] = 8'h06;
DFS[16'h2856] = 8'h0D;
DFS[16'h2857] = 8'h8D;
DFS[16'h2858] = 8'h07;
DFS[16'h2859] = 8'h0D;
DFS[16'h285A] = 8'h8D;
DFS[16'h285B] = 8'h08;
DFS[16'h285C] = 8'h0D;
DFS[16'h285D] = 8'hA9;
DFS[16'h285E] = 8'hFF;
DFS[16'h285F] = 8'h8D;
DFS[16'h2860] = 8'h09;
DFS[16'h2861] = 8'h0D;
DFS[16'h2862] = 8'h8D;
DFS[16'h2863] = 8'h0A;
DFS[16'h2864] = 8'h0D;
DFS[16'h2865] = 8'h8D;
DFS[16'h2866] = 8'h0B;
DFS[16'h2867] = 8'h0D;
DFS[16'h2868] = 8'h4C;
DFS[16'h2869] = 8'h99;
DFS[16'h286A] = 8'hA9;
DFS[16'h286B] = 8'hAD;
DFS[16'h286C] = 8'hFE;
DFS[16'h286D] = 8'h0F;
DFS[16'h286E] = 8'hC9;
DFS[16'h286F] = 8'h55;
DFS[16'h2870] = 8'hD0;
DFS[16'h2871] = 8'h05;
DFS[16'h2872] = 8'hAD;
DFS[16'h2873] = 8'hFF;
DFS[16'h2874] = 8'h0F;
DFS[16'h2875] = 8'hC9;
DFS[16'h2876] = 8'hAA;
DFS[16'h2877] = 8'h60;
DFS[16'h2878] = 8'h4C;
DFS[16'h2879] = 8'hA9;
DFS[16'h287A] = 8'hA9;
DFS[16'h287B] = 8'hAD;
DFS[16'h287C] = 8'hC6;
DFS[16'h287D] = 8'h0F;
DFS[16'h287E] = 8'h0A;
DFS[16'h287F] = 8'h85;
DFS[16'h2880] = 8'hA2;
DFS[16'h2881] = 8'hAD;
DFS[16'h2882] = 8'hC7;
DFS[16'h2883] = 8'h0F;
DFS[16'h2884] = 8'h2A;
DFS[16'h2885] = 8'h85;
DFS[16'h2886] = 8'hA3;
DFS[16'h2887] = 8'hAD;
DFS[16'h2888] = 8'hC8;
DFS[16'h2889] = 8'h0F;
DFS[16'h288A] = 8'h2A;
DFS[16'h288B] = 8'hB0;
DFS[16'h288C] = 8'hEB;
DFS[16'h288D] = 8'h85;
DFS[16'h288E] = 8'hA4;
DFS[16'h288F] = 8'hAD;
DFS[16'h2890] = 8'hC9;
DFS[16'h2891] = 8'h0F;
DFS[16'h2892] = 8'hD0;
DFS[16'h2893] = 8'hE4;
DFS[16'h2894] = 8'h20;
DFS[16'h2895] = 8'h0F;
DFS[16'h2896] = 8'hA6;
DFS[16'h2897] = 8'h20;
DFS[16'h2898] = 8'h6B;
DFS[16'h2899] = 8'hA8;
DFS[16'h289A] = 8'hD0;
DFS[16'h289B] = 8'hDC;
DFS[16'h289C] = 8'hAD;
DFS[16'h289D] = 8'h0B;
DFS[16'h289E] = 8'h0E;
DFS[16'h289F] = 8'hD0;
DFS[16'h28A0] = 8'hD7;
DFS[16'h28A1] = 8'hAD;
DFS[16'h28A2] = 8'h0C;
DFS[16'h28A3] = 8'h0E;
DFS[16'h28A4] = 8'hC9;
DFS[16'h28A5] = 8'h02;
DFS[16'h28A6] = 8'hD0;
DFS[16'h28A7] = 8'hD0;
DFS[16'h28A8] = 8'hAD;
DFS[16'h28A9] = 8'h11;
DFS[16'h28AA] = 8'h0E;
DFS[16'h28AB] = 8'h85;
DFS[16'h28AC] = 8'hA5;
DFS[16'h28AD] = 8'hAD;
DFS[16'h28AE] = 8'h12;
DFS[16'h28AF] = 8'h0E;
DFS[16'h28B0] = 8'h4A;
DFS[16'h28B1] = 8'h66;
DFS[16'h28B2] = 8'hA5;
DFS[16'h28B3] = 8'h4A;
DFS[16'h28B4] = 8'h66;
DFS[16'h28B5] = 8'hA5;
DFS[16'h28B6] = 8'h4A;
DFS[16'h28B7] = 8'h66;
DFS[16'h28B8] = 8'hA5;
DFS[16'h28B9] = 8'h85;
DFS[16'h28BA] = 8'hA6;
DFS[16'h28BB] = 8'hAD;
DFS[16'h28BC] = 8'h0D;
DFS[16'h28BD] = 8'h0E;
DFS[16'h28BE] = 8'h85;
DFS[16'h28BF] = 8'hA7;
DFS[16'h28C0] = 8'hAD;
DFS[16'h28C1] = 8'h0E;
DFS[16'h28C2] = 8'h0E;
DFS[16'h28C3] = 8'h0A;
DFS[16'h28C4] = 8'h2E;
DFS[16'h28C5] = 8'h0F;
DFS[16'h28C6] = 8'h0E;
DFS[16'h28C7] = 8'hB0;
DFS[16'h28C8] = 8'hAF;
DFS[16'h28C9] = 8'h65;
DFS[16'h28CA] = 8'hA2;
DFS[16'h28CB] = 8'h85;
DFS[16'h28CC] = 8'hA2;
DFS[16'h28CD] = 8'hAD;
DFS[16'h28CE] = 8'h0F;
DFS[16'h28CF] = 8'h0E;
DFS[16'h28D0] = 8'h65;
DFS[16'h28D1] = 8'hA3;
DFS[16'h28D2] = 8'h85;
DFS[16'h28D3] = 8'hA3;
DFS[16'h28D4] = 8'h90;
DFS[16'h28D5] = 8'h02;
DFS[16'h28D6] = 8'hE6;
DFS[16'h28D7] = 8'hA4;
DFS[16'h28D8] = 8'h0E;
DFS[16'h28D9] = 8'h16;
DFS[16'h28DA] = 8'h0E;
DFS[16'h28DB] = 8'h2E;
DFS[16'h28DC] = 8'h17;
DFS[16'h28DD] = 8'h0E;
DFS[16'h28DE] = 8'hB0;
DFS[16'h28DF] = 8'h98;
DFS[16'h28E0] = 8'hAE;
DFS[16'h28E1] = 8'h10;
DFS[16'h28E2] = 8'h0E;
DFS[16'h28E3] = 8'h18;
DFS[16'h28E4] = 8'hA5;
DFS[16'h28E5] = 8'hA2;
DFS[16'h28E6] = 8'h6D;
DFS[16'h28E7] = 8'h16;
DFS[16'h28E8] = 8'h0E;
DFS[16'h28E9] = 8'h85;
DFS[16'h28EA] = 8'hA2;
DFS[16'h28EB] = 8'hA5;
DFS[16'h28EC] = 8'hA3;
DFS[16'h28ED] = 8'h6D;
DFS[16'h28EE] = 8'h17;
DFS[16'h28EF] = 8'h0E;
DFS[16'h28F0] = 8'h85;
DFS[16'h28F1] = 8'hA3;
DFS[16'h28F2] = 8'h90;
DFS[16'h28F3] = 8'h02;
DFS[16'h28F4] = 8'hE6;
DFS[16'h28F5] = 8'hA4;
DFS[16'h28F6] = 8'hCA;
DFS[16'h28F7] = 8'hD0;
DFS[16'h28F8] = 8'hEA;
DFS[16'h28F9] = 8'h20;
DFS[16'h28FA] = 8'h0F;
DFS[16'h28FB] = 8'hA6;
DFS[16'h28FC] = 8'hA9;
DFS[16'h28FD] = 8'h00;
DFS[16'h28FE] = 8'h85;
DFS[16'h28FF] = 8'hA8;
DFS[16'h2900] = 8'hA9;
DFS[16'h2901] = 8'h0E;
DFS[16'h2902] = 8'h85;
DFS[16'h2903] = 8'hA9;
DFS[16'h2904] = 8'hA0;
DFS[16'h2905] = 8'h0B;
DFS[16'h2906] = 8'hB1;
DFS[16'h2907] = 8'hA8;
DFS[16'h2908] = 8'h29;
DFS[16'h2909] = 8'h0F;
DFS[16'h290A] = 8'hD0;
DFS[16'h290B] = 8'h10;
DFS[16'h290C] = 8'hA0;
DFS[16'h290D] = 8'h00;
DFS[16'h290E] = 8'hB1;
DFS[16'h290F] = 8'hA8;
DFS[16'h2910] = 8'hD9;
DFS[16'h2911] = 8'hC2;
DFS[16'h2912] = 8'hA9;
DFS[16'h2913] = 8'hD0;
DFS[16'h2914] = 8'h07;
DFS[16'h2915] = 8'hC8;
DFS[16'h2916] = 8'hC0;
DFS[16'h2917] = 8'h0B;
DFS[16'h2918] = 8'hF0;
DFS[16'h2919] = 8'h20;
DFS[16'h291A] = 8'hD0;
DFS[16'h291B] = 8'hF2;
DFS[16'h291C] = 8'h18;
DFS[16'h291D] = 8'hA5;
DFS[16'h291E] = 8'hA8;
DFS[16'h291F] = 8'h69;
DFS[16'h2920] = 8'h20;
DFS[16'h2921] = 8'h85;
DFS[16'h2922] = 8'hA8;
DFS[16'h2923] = 8'hD0;
DFS[16'h2924] = 8'hDF;
DFS[16'h2925] = 8'h20;
DFS[16'h2926] = 8'h00;
DFS[16'h2927] = 8'hA0;
DFS[16'h2928] = 8'hFF;
DFS[16'h2929] = 8'h49;
DFS[16'h292A] = 8'h6D;
DFS[16'h292B] = 8'h61;
DFS[16'h292C] = 8'h67;
DFS[16'h292D] = 8'h65;
DFS[16'h292E] = 8'h20;
DFS[16'h292F] = 8'h6E;
DFS[16'h2930] = 8'h6F;
DFS[16'h2931] = 8'h74;
DFS[16'h2932] = 8'h20;
DFS[16'h2933] = 8'h66;
DFS[16'h2934] = 8'h6F;
DFS[16'h2935] = 8'h75;
DFS[16'h2936] = 8'h6E;
DFS[16'h2937] = 8'h64;
DFS[16'h2938] = 8'h21;
DFS[16'h2939] = 8'h00;
DFS[16'h293A] = 8'h18;
DFS[16'h293B] = 8'hA5;
DFS[16'h293C] = 8'hA2;
DFS[16'h293D] = 8'h65;
DFS[16'h293E] = 8'hA5;
DFS[16'h293F] = 8'h85;
DFS[16'h2940] = 8'hA2;
DFS[16'h2941] = 8'hA5;
DFS[16'h2942] = 8'hA3;
DFS[16'h2943] = 8'h65;
DFS[16'h2944] = 8'hA6;
DFS[16'h2945] = 8'h85;
DFS[16'h2946] = 8'hA3;
DFS[16'h2947] = 8'h90;
DFS[16'h2948] = 8'h02;
DFS[16'h2949] = 8'hE6;
DFS[16'h294A] = 8'hA4;
DFS[16'h294B] = 8'hA0;
DFS[16'h294C] = 8'h1B;
DFS[16'h294D] = 8'hB1;
DFS[16'h294E] = 8'hA8;
DFS[16'h294F] = 8'h48;
DFS[16'h2950] = 8'h88;
DFS[16'h2951] = 8'hB1;
DFS[16'h2952] = 8'hA8;
DFS[16'h2953] = 8'h38;
DFS[16'h2954] = 8'hE9;
DFS[16'h2955] = 8'h02;
DFS[16'h2956] = 8'h85;
DFS[16'h2957] = 8'hA8;
DFS[16'h2958] = 8'h68;
DFS[16'h2959] = 8'hE9;
DFS[16'h295A] = 8'h00;
DFS[16'h295B] = 8'h85;
DFS[16'h295C] = 8'hA9;
DFS[16'h295D] = 8'h05;
DFS[16'h295E] = 8'hA8;
DFS[16'h295F] = 8'hF0;
DFS[16'h2960] = 8'h1A;
DFS[16'h2961] = 8'h06;
DFS[16'h2962] = 8'hA8;
DFS[16'h2963] = 8'h26;
DFS[16'h2964] = 8'hA9;
DFS[16'h2965] = 8'hA6;
DFS[16'h2966] = 8'hA7;
DFS[16'h2967] = 8'h18;
DFS[16'h2968] = 8'hA5;
DFS[16'h2969] = 8'hA2;
DFS[16'h296A] = 8'h65;
DFS[16'h296B] = 8'hA8;
DFS[16'h296C] = 8'h85;
DFS[16'h296D] = 8'hA2;
DFS[16'h296E] = 8'hA5;
DFS[16'h296F] = 8'hA3;
DFS[16'h2970] = 8'h65;
DFS[16'h2971] = 8'hA9;
DFS[16'h2972] = 8'h85;
DFS[16'h2973] = 8'hA3;
DFS[16'h2974] = 8'h90;
DFS[16'h2975] = 8'h02;
DFS[16'h2976] = 8'hE6;
DFS[16'h2977] = 8'hA4;
DFS[16'h2978] = 8'hCA;
DFS[16'h2979] = 8'hD0;
DFS[16'h297A] = 8'hEC;
DFS[16'h297B] = 8'hA5;
DFS[16'h297C] = 8'hA2;
DFS[16'h297D] = 8'h8D;
DFS[16'h297E] = 8'h06;
DFS[16'h297F] = 8'h0D;
DFS[16'h2980] = 8'h49;
DFS[16'h2981] = 8'hFF;
DFS[16'h2982] = 8'h8D;
DFS[16'h2983] = 8'h09;
DFS[16'h2984] = 8'h0D;
DFS[16'h2985] = 8'hA5;
DFS[16'h2986] = 8'hA3;
DFS[16'h2987] = 8'h8D;
DFS[16'h2988] = 8'h07;
DFS[16'h2989] = 8'h0D;
DFS[16'h298A] = 8'h49;
DFS[16'h298B] = 8'hFF;
DFS[16'h298C] = 8'h8D;
DFS[16'h298D] = 8'h0A;
DFS[16'h298E] = 8'h0D;
DFS[16'h298F] = 8'hA5;
DFS[16'h2990] = 8'hA4;
DFS[16'h2991] = 8'h8D;
DFS[16'h2992] = 8'h08;
DFS[16'h2993] = 8'h0D;
DFS[16'h2994] = 8'h49;
DFS[16'h2995] = 8'hFF;
DFS[16'h2996] = 8'h8D;
DFS[16'h2997] = 8'h0B;
DFS[16'h2998] = 8'h0D;
DFS[16'h2999] = 8'hA9;
DFS[16'h299A] = 8'h54;
DFS[16'h299B] = 8'h8D;
DFS[16'h299C] = 8'h05;
DFS[16'h299D] = 8'h0D;
DFS[16'h299E] = 8'hA2;
DFS[16'h299F] = 8'h00;
DFS[16'h29A0] = 8'h68;
DFS[16'h29A1] = 8'h95;
DFS[16'h29A2] = 8'hA2;
DFS[16'h29A3] = 8'hE8;
DFS[16'h29A4] = 8'hE0;
DFS[16'h29A5] = 8'h08;
DFS[16'h29A6] = 8'hD0;
DFS[16'h29A7] = 8'hF8;
DFS[16'h29A8] = 8'h60;
DFS[16'h29A9] = 8'h20;
DFS[16'h29AA] = 8'h00;
DFS[16'h29AB] = 8'hA0;
DFS[16'h29AC] = 8'hFF;
DFS[16'h29AD] = 8'h55;
DFS[16'h29AE] = 8'h6E;
DFS[16'h29AF] = 8'h72;
DFS[16'h29B0] = 8'h65;
DFS[16'h29B1] = 8'h63;
DFS[16'h29B2] = 8'h6F;
DFS[16'h29B3] = 8'h67;
DFS[16'h29B4] = 8'h6E;
DFS[16'h29B5] = 8'h69;
DFS[16'h29B6] = 8'h73;
DFS[16'h29B7] = 8'h65;
DFS[16'h29B8] = 8'h64;
DFS[16'h29B9] = 8'h20;
DFS[16'h29BA] = 8'h66;
DFS[16'h29BB] = 8'h6F;
DFS[16'h29BC] = 8'h72;
DFS[16'h29BD] = 8'h6D;
DFS[16'h29BE] = 8'h61;
DFS[16'h29BF] = 8'h74;
DFS[16'h29C0] = 8'h21;
DFS[16'h29C1] = 8'h00;
DFS[16'h29C2] = 8'h42;
DFS[16'h29C3] = 8'h45;
DFS[16'h29C4] = 8'h45;
DFS[16'h29C5] = 8'h42;
DFS[16'h29C6] = 8'h20;
DFS[16'h29C7] = 8'h20;
DFS[16'h29C8] = 8'h20;
DFS[16'h29C9] = 8'h20;
DFS[16'h29CA] = 8'h4D;
DFS[16'h29CB] = 8'h4D;
DFS[16'h29CC] = 8'h42;
DFS[16'h29CD] = 8'h08;
DFS[16'h29CE] = 8'hAA;
DFS[16'h29CF] = 8'h20;
DFS[16'h29D0] = 8'h02;
DFS[16'h29D1] = 8'hAA;
DFS[16'h29D2] = 8'h85;
DFS[16'h29D3] = 8'hB2;
DFS[16'h29D4] = 8'h48;
DFS[16'h29D5] = 8'h20;
DFS[16'h29D6] = 8'h1E;
DFS[16'h29D7] = 8'hAA;
DFS[16'h29D8] = 8'h8A;
DFS[16'h29D9] = 8'hE5;
DFS[16'h29DA] = 8'hB0;
DFS[16'h29DB] = 8'hAA;
DFS[16'h29DC] = 8'h68;
DFS[16'h29DD] = 8'h20;
DFS[16'h29DE] = 8'h02;
DFS[16'h29DF] = 8'hAA;
DFS[16'h29E0] = 8'h48;
DFS[16'h29E1] = 8'h20;
DFS[16'h29E2] = 8'h1E;
DFS[16'h29E3] = 8'hAA;
DFS[16'h29E4] = 8'hA5;
DFS[16'h29E5] = 8'hB2;
DFS[16'h29E6] = 8'hE5;
DFS[16'h29E7] = 8'hB0;
DFS[16'h29E8] = 8'h0A;
DFS[16'h29E9] = 8'h0A;
DFS[16'h29EA] = 8'h0A;
DFS[16'h29EB] = 8'h0A;
DFS[16'h29EC] = 8'h85;
DFS[16'h29ED] = 8'hB2;
DFS[16'h29EE] = 8'h8A;
DFS[16'h29EF] = 8'h05;
DFS[16'h29F0] = 8'hB2;
DFS[16'h29F1] = 8'hAA;
DFS[16'h29F2] = 8'h68;
DFS[16'h29F3] = 8'h28;
DFS[16'h29F4] = 8'h90;
DFS[16'h29F5] = 8'h0B;
DFS[16'h29F6] = 8'h48;
DFS[16'h29F7] = 8'h8A;
DFS[16'h29F8] = 8'hF8;
DFS[16'h29F9] = 8'h18;
DFS[16'h29FA] = 8'h69;
DFS[16'h29FB] = 8'h56;
DFS[16'h29FC] = 8'hAA;
DFS[16'h29FD] = 8'h68;
DFS[16'h29FE] = 8'h69;
DFS[16'h29FF] = 8'h02;
DFS[16'h2A00] = 8'hD8;
DFS[16'h2A01] = 8'h60;
DFS[16'h2A02] = 8'hA0;
DFS[16'h2A03] = 8'h00;
DFS[16'h2A04] = 8'h84;
DFS[16'h2A05] = 8'hB1;
DFS[16'h2A06] = 8'hA0;
DFS[16'h2A07] = 8'hA0;
DFS[16'h2A08] = 8'h84;
DFS[16'h2A09] = 8'hB0;
DFS[16'h2A0A] = 8'hA0;
DFS[16'h2A0B] = 8'h05;
DFS[16'h2A0C] = 8'hC5;
DFS[16'h2A0D] = 8'hB0;
DFS[16'h2A0E] = 8'h90;
DFS[16'h2A0F] = 8'h04;
DFS[16'h2A10] = 8'h38;
DFS[16'h2A11] = 8'hE5;
DFS[16'h2A12] = 8'hB0;
DFS[16'h2A13] = 8'h38;
DFS[16'h2A14] = 8'h26;
DFS[16'h2A15] = 8'hB1;
DFS[16'h2A16] = 8'h46;
DFS[16'h2A17] = 8'hB0;
DFS[16'h2A18] = 8'h88;
DFS[16'h2A19] = 8'hD0;
DFS[16'h2A1A] = 8'hF1;
DFS[16'h2A1B] = 8'hA5;
DFS[16'h2A1C] = 8'hB1;
DFS[16'h2A1D] = 8'h60;
DFS[16'h2A1E] = 8'h48;
DFS[16'h2A1F] = 8'h0A;
DFS[16'h2A20] = 8'h0A;
DFS[16'h2A21] = 8'h0A;
DFS[16'h2A22] = 8'h85;
DFS[16'h2A23] = 8'hB0;
DFS[16'h2A24] = 8'h68;
DFS[16'h2A25] = 8'h0A;
DFS[16'h2A26] = 8'h18;
DFS[16'h2A27] = 8'h65;
DFS[16'h2A28] = 8'hB0;
DFS[16'h2A29] = 8'h85;
DFS[16'h2A2A] = 8'hB0;
DFS[16'h2A2B] = 8'h38;
DFS[16'h2A2C] = 8'h60;
DFS[16'h2A2D] = 8'hE0;
DFS[16'h2A2E] = 8'hFF;
DFS[16'h2A2F] = 8'hF0;
DFS[16'h2A30] = 8'h35;
DFS[16'h2A31] = 8'hBD;
DFS[16'h2A32] = 8'h10;
DFS[16'h2A33] = 8'h0D;
DFS[16'h2A34] = 8'h30;
DFS[16'h2A35] = 8'h30;
DFS[16'h2A36] = 8'h49;
DFS[16'h2A37] = 8'hFF;
DFS[16'h2A38] = 8'hDD;
DFS[16'h2A39] = 8'h18;
DFS[16'h2A3A] = 8'h0D;
DFS[16'h2A3B] = 8'hD0;
DFS[16'h2A3C] = 8'h24;
DFS[16'h2A3D] = 8'hBD;
DFS[16'h2A3E] = 8'h0C;
DFS[16'h2A3F] = 8'h0D;
DFS[16'h2A40] = 8'h49;
DFS[16'h2A41] = 8'hFF;
DFS[16'h2A42] = 8'hDD;
DFS[16'h2A43] = 8'h14;
DFS[16'h2A44] = 8'h0D;
DFS[16'h2A45] = 8'hD0;
DFS[16'h2A46] = 8'h1A;
DFS[16'h2A47] = 8'hBD;
DFS[16'h2A48] = 8'h1C;
DFS[16'h2A49] = 8'h0D;
DFS[16'h2A4A] = 8'hC9;
DFS[16'h2A4B] = 8'h54;
DFS[16'h2A4C] = 8'hF0;
DFS[16'h2A4D] = 8'h29;
DFS[16'h2A4E] = 8'h20;
DFS[16'h2A4F] = 8'h00;
DFS[16'h2A50] = 8'hA0;
DFS[16'h2A51] = 8'hC9;
DFS[16'h2A52] = 8'h44;
DFS[16'h2A53] = 8'h69;
DFS[16'h2A54] = 8'h73;
DFS[16'h2A55] = 8'h6B;
DFS[16'h2A56] = 8'h20;
DFS[16'h2A57] = 8'h72;
DFS[16'h2A58] = 8'h65;
DFS[16'h2A59] = 8'h61;
DFS[16'h2A5A] = 8'h64;
DFS[16'h2A5B] = 8'h20;
DFS[16'h2A5C] = 8'h6F;
DFS[16'h2A5D] = 8'h6E;
DFS[16'h2A5E] = 8'h6C;
DFS[16'h2A5F] = 8'h79;
DFS[16'h2A60] = 8'h00;
DFS[16'h2A61] = 8'hA9;
DFS[16'h2A62] = 8'hFF;
DFS[16'h2A63] = 8'h9D;
DFS[16'h2A64] = 8'h10;
DFS[16'h2A65] = 8'h0D;
DFS[16'h2A66] = 8'h20;
DFS[16'h2A67] = 8'h00;
DFS[16'h2A68] = 8'hA0;
DFS[16'h2A69] = 8'hC7;
DFS[16'h2A6A] = 8'h4E;
DFS[16'h2A6B] = 8'h6F;
DFS[16'h2A6C] = 8'h20;
DFS[16'h2A6D] = 8'h64;
DFS[16'h2A6E] = 8'h69;
DFS[16'h2A6F] = 8'h73;
DFS[16'h2A70] = 8'h6B;
DFS[16'h2A71] = 8'h00;
DFS[16'h2A72] = 8'hA9;
DFS[16'h2A73] = 8'h54;
DFS[16'h2A74] = 8'h9D;
DFS[16'h2A75] = 8'h1C;
DFS[16'h2A76] = 8'h0D;
DFS[16'h2A77] = 8'h60;
DFS[16'h2A78] = 8'hA9;
DFS[16'h2A79] = 8'h00;
DFS[16'h2A7A] = 8'h9D;
DFS[16'h2A7B] = 8'h1C;
DFS[16'h2A7C] = 8'h0D;
DFS[16'h2A7D] = 8'h60;
DFS[16'h2A7E] = 8'hBD;
DFS[16'h2A7F] = 8'h10;
DFS[16'h2A80] = 8'h0D;
DFS[16'h2A81] = 8'h30;
DFS[16'h2A82] = 8'hE3;
DFS[16'h2A83] = 8'h6A;
DFS[16'h2A84] = 8'hBD;
DFS[16'h2A85] = 8'h0C;
DFS[16'h2A86] = 8'h0D;
DFS[16'h2A87] = 8'h08;
DFS[16'h2A88] = 8'hAA;
DFS[16'h2A89] = 8'hA9;
DFS[16'h2A8A] = 8'h00;
DFS[16'h2A8B] = 8'h85;
DFS[16'h2A8C] = 8'hA2;
DFS[16'h2A8D] = 8'h2A;
DFS[16'h2A8E] = 8'h48;
DFS[16'h2A8F] = 8'h85;
DFS[16'h2A90] = 8'hA4;
DFS[16'h2A91] = 8'h8A;
DFS[16'h2A92] = 8'h0A;
DFS[16'h2A93] = 8'h26;
DFS[16'h2A94] = 8'hA4;
DFS[16'h2A95] = 8'h85;
DFS[16'h2A96] = 8'hA3;
DFS[16'h2A97] = 8'h8A;
DFS[16'h2A98] = 8'h65;
DFS[16'h2A99] = 8'hA3;
DFS[16'h2A9A] = 8'h85;
DFS[16'h2A9B] = 8'hA3;
DFS[16'h2A9C] = 8'h68;
DFS[16'h2A9D] = 8'h69;
DFS[16'h2A9E] = 8'h00;
DFS[16'h2A9F] = 8'h65;
DFS[16'h2AA0] = 8'hA4;
DFS[16'h2AA1] = 8'h85;
DFS[16'h2AA2] = 8'hA4;
DFS[16'h2AA3] = 8'h66;
DFS[16'h2AA4] = 8'hA2;
DFS[16'h2AA5] = 8'h8A;
DFS[16'h2AA6] = 8'h28;
DFS[16'h2AA7] = 8'h6A;
DFS[16'h2AA8] = 8'h66;
DFS[16'h2AA9] = 8'hA2;
DFS[16'h2AAA] = 8'h4A;
DFS[16'h2AAB] = 8'h66;
DFS[16'h2AAC] = 8'hA2;
DFS[16'h2AAD] = 8'h4A;
DFS[16'h2AAE] = 8'h66;
DFS[16'h2AAF] = 8'hA2;
DFS[16'h2AB0] = 8'h65;
DFS[16'h2AB1] = 8'hA3;
DFS[16'h2AB2] = 8'h85;
DFS[16'h2AB3] = 8'hA3;
DFS[16'h2AB4] = 8'hA5;
DFS[16'h2AB5] = 8'hA4;
DFS[16'h2AB6] = 8'h69;
DFS[16'h2AB7] = 8'h00;
DFS[16'h2AB8] = 8'h85;
DFS[16'h2AB9] = 8'hA4;
DFS[16'h2ABA] = 8'h20;
DFS[16'h2ABB] = 8'h17;
DFS[16'h2ABC] = 8'hA8;
DFS[16'h2ABD] = 8'h38;
DFS[16'h2ABE] = 8'hA5;
DFS[16'h2ABF] = 8'hA2;
DFS[16'h2AC0] = 8'h09;
DFS[16'h2AC1] = 8'h1F;
DFS[16'h2AC2] = 8'h6D;
DFS[16'h2AC3] = 8'h06;
DFS[16'h2AC4] = 8'h0D;
DFS[16'h2AC5] = 8'h85;
DFS[16'h2AC6] = 8'hA2;
DFS[16'h2AC7] = 8'hA5;
DFS[16'h2AC8] = 8'hA3;
DFS[16'h2AC9] = 8'h6D;
DFS[16'h2ACA] = 8'h07;
DFS[16'h2ACB] = 8'h0D;
DFS[16'h2ACC] = 8'h85;
DFS[16'h2ACD] = 8'hA3;
DFS[16'h2ACE] = 8'hA5;
DFS[16'h2ACF] = 8'hA4;
DFS[16'h2AD0] = 8'h6D;
DFS[16'h2AD1] = 8'h08;
DFS[16'h2AD2] = 8'h0D;
DFS[16'h2AD3] = 8'h85;
DFS[16'h2AD4] = 8'hA4;
DFS[16'h2AD5] = 8'h60;
DFS[16'h2AD6] = 8'hA5;
DFS[16'h2AD7] = 8'hBE;
DFS[16'h2AD8] = 8'h85;
DFS[16'h2AD9] = 8'hA0;
DFS[16'h2ADA] = 8'hA5;
DFS[16'h2ADB] = 8'hBF;
DFS[16'h2ADC] = 8'h85;
DFS[16'h2ADD] = 8'hA1;
DFS[16'h2ADE] = 8'hA6;
DFS[16'h2ADF] = 8'hCF;
DFS[16'h2AE0] = 8'h20;
DFS[16'h2AE1] = 8'h7E;
DFS[16'h2AE2] = 8'hAA;
DFS[16'h2AE3] = 8'h18;
DFS[16'h2AE4] = 8'hA5;
DFS[16'h2AE5] = 8'hC5;
DFS[16'h2AE6] = 8'h65;
DFS[16'h2AE7] = 8'hA2;
DFS[16'h2AE8] = 8'h85;
DFS[16'h2AE9] = 8'hA2;
DFS[16'h2AEA] = 8'hA5;
DFS[16'h2AEB] = 8'hC4;
DFS[16'h2AEC] = 8'h29;
DFS[16'h2AED] = 8'h03;
DFS[16'h2AEE] = 8'h48;
DFS[16'h2AEF] = 8'h65;
DFS[16'h2AF0] = 8'hA3;
DFS[16'h2AF1] = 8'h85;
DFS[16'h2AF2] = 8'hA3;
DFS[16'h2AF3] = 8'h90;
DFS[16'h2AF4] = 8'h02;
DFS[16'h2AF5] = 8'hE6;
DFS[16'h2AF6] = 8'hA4;
DFS[16'h2AF7] = 8'hA5;
DFS[16'h2AF8] = 8'hC3;
DFS[16'h2AF9] = 8'h85;
DFS[16'h2AFA] = 8'hA5;
DFS[16'h2AFB] = 8'hA5;
DFS[16'h2AFC] = 8'hC4;
DFS[16'h2AFD] = 8'h4A;
DFS[16'h2AFE] = 8'h4A;
DFS[16'h2AFF] = 8'h4A;
DFS[16'h2B00] = 8'h4A;
DFS[16'h2B01] = 8'h29;
DFS[16'h2B02] = 8'h03;
DFS[16'h2B03] = 8'hD0;
DFS[16'h2B04] = 8'h1E;
DFS[16'h2B05] = 8'hA5;
DFS[16'h2B06] = 8'hC2;
DFS[16'h2B07] = 8'h85;
DFS[16'h2B08] = 8'hA7;
DFS[16'h2B09] = 8'hF0;
DFS[16'h2B0A] = 8'h04;
DFS[16'h2B0B] = 8'hE6;
DFS[16'h2B0C] = 8'hA5;
DFS[16'h2B0D] = 8'hF0;
DFS[16'h2B0E] = 8'h14;
DFS[16'h2B0F] = 8'h18;
DFS[16'h2B10] = 8'hA5;
DFS[16'h2B11] = 8'hC5;
DFS[16'h2B12] = 8'h65;
DFS[16'h2B13] = 8'hA5;
DFS[16'h2B14] = 8'hAA;
DFS[16'h2B15] = 8'h68;
DFS[16'h2B16] = 8'h69;
DFS[16'h2B17] = 8'h00;
DFS[16'h2B18] = 8'hC9;
DFS[16'h2B19] = 8'h03;
DFS[16'h2B1A] = 8'h90;
DFS[16'h2B1B] = 8'h06;
DFS[16'h2B1C] = 8'hD0;
DFS[16'h2B1D] = 8'h17;
DFS[16'h2B1E] = 8'hE0;
DFS[16'h2B1F] = 8'h21;
DFS[16'h2B20] = 8'hB0;
DFS[16'h2B21] = 8'h13;
DFS[16'h2B22] = 8'h60;
DFS[16'h2B23] = 8'h20;
DFS[16'h2B24] = 8'h00;
DFS[16'h2B25] = 8'hA0;
DFS[16'h2B26] = 8'hFF;
DFS[16'h2B27] = 8'h42;
DFS[16'h2B28] = 8'h6C;
DFS[16'h2B29] = 8'h6F;
DFS[16'h2B2A] = 8'h63;
DFS[16'h2B2B] = 8'h6B;
DFS[16'h2B2C] = 8'h20;
DFS[16'h2B2D] = 8'h74;
DFS[16'h2B2E] = 8'h6F;
DFS[16'h2B2F] = 8'h6F;
DFS[16'h2B30] = 8'h20;
DFS[16'h2B31] = 8'h62;
DFS[16'h2B32] = 8'h69;
DFS[16'h2B33] = 8'h67;
DFS[16'h2B34] = 8'h00;
DFS[16'h2B35] = 8'h20;
DFS[16'h2B36] = 8'h00;
DFS[16'h2B37] = 8'hA0;
DFS[16'h2B38] = 8'hFF;
DFS[16'h2B39] = 8'h44;
DFS[16'h2B3A] = 8'h69;
DFS[16'h2B3B] = 8'h73;
DFS[16'h2B3C] = 8'h6B;
DFS[16'h2B3D] = 8'h20;
DFS[16'h2B3E] = 8'h6F;
DFS[16'h2B3F] = 8'h76;
DFS[16'h2B40] = 8'h65;
DFS[16'h2B41] = 8'h72;
DFS[16'h2B42] = 8'h66;
DFS[16'h2B43] = 8'h6C;
DFS[16'h2B44] = 8'h6F;
DFS[16'h2B45] = 8'h77;
DFS[16'h2B46] = 8'h00;
DFS[16'h2B47] = 8'h20;
DFS[16'h2B48] = 8'h4D;
DFS[16'h2B49] = 8'h83;
DFS[16'h2B4A] = 8'h20;
DFS[16'h2B4B] = 8'h58;
DFS[16'h2B4C] = 8'h83;
DFS[16'h2B4D] = 8'h20;
DFS[16'h2B4E] = 8'hEC;
DFS[16'h2B4F] = 8'hA4;
DFS[16'h2B50] = 8'hA6;
DFS[16'h2B51] = 8'hCF;
DFS[16'h2B52] = 8'h8E;
DFS[16'h2B53] = 8'h20;
DFS[16'h2B54] = 8'h0D;
DFS[16'h2B55] = 8'h20;
DFS[16'h2B56] = 8'h7E;
DFS[16'h2B57] = 8'hAA;
DFS[16'h2B58] = 8'h20;
DFS[16'h2B59] = 8'h0F;
DFS[16'h2B5A] = 8'hA6;
DFS[16'h2B5B] = 8'hA5;
DFS[16'h2B5C] = 8'hCF;
DFS[16'h2B5D] = 8'h8D;
DFS[16'h2B5E] = 8'h82;
DFS[16'h2B5F] = 8'h10;
DFS[16'h2B60] = 8'h60;
DFS[16'h2B61] = 8'h20;
DFS[16'h2B62] = 8'hEC;
DFS[16'h2B63] = 8'hA4;
DFS[16'h2B64] = 8'hA6;
DFS[16'h2B65] = 8'hCF;
DFS[16'h2B66] = 8'h20;
DFS[16'h2B67] = 8'h2D;
DFS[16'h2B68] = 8'hAA;
DFS[16'h2B69] = 8'h20;
DFS[16'h2B6A] = 8'h7E;
DFS[16'h2B6B] = 8'hAA;
DFS[16'h2B6C] = 8'h4C;
DFS[16'h2B6D] = 8'h28;
DFS[16'h2B6E] = 8'hA6;
DFS[16'h2B6F] = 8'h08;
DFS[16'h2B70] = 8'h48;
DFS[16'h2B71] = 8'hA0;
DFS[16'h2B72] = 8'hFF;
DFS[16'h2B73] = 8'h8C;
DFS[16'h2B74] = 8'h82;
DFS[16'h2B75] = 8'h10;
DFS[16'h2B76] = 8'hC8;
DFS[16'h2B77] = 8'h98;
DFS[16'h2B78] = 8'h99;
DFS[16'h2B79] = 8'h00;
DFS[16'h2B7A] = 8'h0E;
DFS[16'h2B7B] = 8'h99;
DFS[16'h2B7C] = 8'h00;
DFS[16'h2B7D] = 8'h0F;
DFS[16'h2B7E] = 8'hC8;
DFS[16'h2B7F] = 8'hD0;
DFS[16'h2B80] = 8'hF7;
DFS[16'h2B81] = 8'hA9;
DFS[16'h2B82] = 8'h03;
DFS[16'h2B83] = 8'h8D;
DFS[16'h2B84] = 8'h06;
DFS[16'h2B85] = 8'h0F;
DFS[16'h2B86] = 8'hA9;
DFS[16'h2B87] = 8'h20;
DFS[16'h2B88] = 8'h8D;
DFS[16'h2B89] = 8'h07;
DFS[16'h2B8A] = 8'h0F;
DFS[16'h2B8B] = 8'h20;
DFS[16'h2B8C] = 8'hEC;
DFS[16'h2B8D] = 8'hA4;
DFS[16'h2B8E] = 8'h68;
DFS[16'h2B8F] = 8'h28;
DFS[16'h2B90] = 8'h20;
DFS[16'h2B91] = 8'h87;
DFS[16'h2B92] = 8'hAA;
DFS[16'h2B93] = 8'h4C;
DFS[16'h2B94] = 8'h28;
DFS[16'h2B95] = 8'hA6;
DFS[16'h2B96] = 8'h20;
DFS[16'h2B97] = 8'hEC;
DFS[16'h2B98] = 8'hA4;
DFS[16'h2B99] = 8'h20;
DFS[16'h2B9A] = 8'hD6;
DFS[16'h2B9B] = 8'hAA;
DFS[16'h2B9C] = 8'h20;
DFS[16'h2B9D] = 8'h42;
DFS[16'h2B9E] = 8'hA6;
DFS[16'h2B9F] = 8'h20;
DFS[16'h2BA0] = 8'hCD;
DFS[16'h2BA1] = 8'hA0;
DFS[16'h2BA2] = 8'hA9;
DFS[16'h2BA3] = 8'h01;
DFS[16'h2BA4] = 8'h60;
DFS[16'h2BA5] = 8'h20;
DFS[16'h2BA6] = 8'hEC;
DFS[16'h2BA7] = 8'hA4;
DFS[16'h2BA8] = 8'h20;
DFS[16'h2BA9] = 8'hD6;
DFS[16'h2BAA] = 8'hAA;
DFS[16'h2BAB] = 8'hA6;
DFS[16'h2BAC] = 8'hCF;
DFS[16'h2BAD] = 8'h20;
DFS[16'h2BAE] = 8'h2D;
DFS[16'h2BAF] = 8'hAA;
DFS[16'h2BB0] = 8'h20;
DFS[16'h2BB1] = 8'hEF;
DFS[16'h2BB2] = 8'hA6;
DFS[16'h2BB3] = 8'h20;
DFS[16'h2BB4] = 8'hCD;
DFS[16'h2BB5] = 8'hA0;
DFS[16'h2BB6] = 8'hA9;
DFS[16'h2BB7] = 8'h01;
DFS[16'h2BB8] = 8'h60;
DFS[16'h2BB9] = 8'hA8;
DFS[16'h2BBA] = 8'hC8;
DFS[16'h2BBB] = 8'h98;
DFS[16'h2BBC] = 8'hD0;
DFS[16'h2BBD] = 8'h01;
DFS[16'h2BBE] = 8'h38;
DFS[16'h2BBF] = 8'h2A;
DFS[16'h2BC0] = 8'h2A;
DFS[16'h2BC1] = 8'h2A;
DFS[16'h2BC2] = 8'h2A;
DFS[16'h2BC3] = 8'h2A;
DFS[16'h2BC4] = 8'h48;
DFS[16'h2BC5] = 8'h29;
DFS[16'h2BC6] = 8'h1F;
DFS[16'h2BC7] = 8'hA8;
DFS[16'h2BC8] = 8'h68;
DFS[16'h2BC9] = 8'h09;
DFS[16'h2BCA] = 8'h1F;
DFS[16'h2BCB] = 8'h6A;
DFS[16'h2BCC] = 8'h60;
DFS[16'h2BCD] = 8'h20;
DFS[16'h2BCE] = 8'hB9;
DFS[16'h2BCF] = 8'hAB;
DFS[16'h2BD0] = 8'h48;
DFS[16'h2BD1] = 8'h8A;
DFS[16'h2BD2] = 8'h48;
DFS[16'h2BD3] = 8'h98;
DFS[16'h2BD4] = 8'h48;
DFS[16'h2BD5] = 8'h20;
DFS[16'h2BD6] = 8'h98;
DFS[16'h2BD7] = 8'hAC;
DFS[16'h2BD8] = 8'h68;
DFS[16'h2BD9] = 8'h6A;
DFS[16'h2BDA] = 8'h68;
DFS[16'h2BDB] = 8'hAA;
DFS[16'h2BDC] = 8'h68;
DFS[16'h2BDD] = 8'hA8;
DFS[16'h2BDE] = 8'hB0;
DFS[16'h2BDF] = 8'h04;
DFS[16'h2BE0] = 8'hB9;
DFS[16'h2BE1] = 8'h00;
DFS[16'h2BE2] = 8'h0E;
DFS[16'h2BE3] = 8'h60;
DFS[16'h2BE4] = 8'hB9;
DFS[16'h2BE5] = 8'h00;
DFS[16'h2BE6] = 8'h0F;
DFS[16'h2BE7] = 8'h60;
DFS[16'h2BE8] = 8'h08;
DFS[16'h2BE9] = 8'h48;
DFS[16'h2BEA] = 8'h8D;
DFS[16'h2BEB] = 8'h5F;
DFS[16'h2BEC] = 8'h0D;
DFS[16'h2BED] = 8'hA9;
DFS[16'h2BEE] = 8'h00;
DFS[16'h2BEF] = 8'h2A;
DFS[16'h2BF0] = 8'h8D;
DFS[16'h2BF1] = 8'h60;
DFS[16'h2BF2] = 8'h0D;
DFS[16'h2BF3] = 8'h8E;
DFS[16'h2BF4] = 8'h61;
DFS[16'h2BF5] = 8'h0D;
DFS[16'h2BF6] = 8'hA2;
DFS[16'h2BF7] = 8'h03;
DFS[16'h2BF8] = 8'hEC;
DFS[16'h2BF9] = 8'h61;
DFS[16'h2BFA] = 8'h0D;
DFS[16'h2BFB] = 8'hF0;
DFS[16'h2BFC] = 8'h15;
DFS[16'h2BFD] = 8'hBD;
DFS[16'h2BFE] = 8'h0C;
DFS[16'h2BFF] = 8'h0D;
DFS[16'h2C00] = 8'hCD;
DFS[16'h2C01] = 8'h5F;
DFS[16'h2C02] = 8'h0D;
DFS[16'h2C03] = 8'hD0;
DFS[16'h2C04] = 8'h0D;
DFS[16'h2C05] = 8'hBD;
DFS[16'h2C06] = 8'h10;
DFS[16'h2C07] = 8'h0D;
DFS[16'h2C08] = 8'hCD;
DFS[16'h2C09] = 8'h60;
DFS[16'h2C0A] = 8'h0D;
DFS[16'h2C0B] = 8'hD0;
DFS[16'h2C0C] = 8'h05;
DFS[16'h2C0D] = 8'hA9;
DFS[16'h2C0E] = 8'hFF;
DFS[16'h2C0F] = 8'h9D;
DFS[16'h2C10] = 8'h10;
DFS[16'h2C11] = 8'h0D;
DFS[16'h2C12] = 8'hCA;
DFS[16'h2C13] = 8'h10;
DFS[16'h2C14] = 8'hE3;
DFS[16'h2C15] = 8'hAE;
DFS[16'h2C16] = 8'h61;
DFS[16'h2C17] = 8'h0D;
DFS[16'h2C18] = 8'h68;
DFS[16'h2C19] = 8'h28;
DFS[16'h2C1A] = 8'h60;
DFS[16'h2C1B] = 8'h08;
DFS[16'h2C1C] = 8'h48;
DFS[16'h2C1D] = 8'h9D;
DFS[16'h2C1E] = 8'h0C;
DFS[16'h2C1F] = 8'h0D;
DFS[16'h2C20] = 8'h49;
DFS[16'h2C21] = 8'hFF;
DFS[16'h2C22] = 8'h9D;
DFS[16'h2C23] = 8'h14;
DFS[16'h2C24] = 8'h0D;
DFS[16'h2C25] = 8'hA9;
DFS[16'h2C26] = 8'h00;
DFS[16'h2C27] = 8'h2A;
DFS[16'h2C28] = 8'h9D;
DFS[16'h2C29] = 8'h10;
DFS[16'h2C2A] = 8'h0D;
DFS[16'h2C2B] = 8'h49;
DFS[16'h2C2C] = 8'hFF;
DFS[16'h2C2D] = 8'h9D;
DFS[16'h2C2E] = 8'h18;
DFS[16'h2C2F] = 8'h0D;
DFS[16'h2C30] = 8'h68;
DFS[16'h2C31] = 8'h28;
DFS[16'h2C32] = 8'h20;
DFS[16'h2C33] = 8'hE8;
DFS[16'h2C34] = 8'hAB;
DFS[16'h2C35] = 8'h20;
DFS[16'h2C36] = 8'hCD;
DFS[16'h2C37] = 8'hAB;
DFS[16'h2C38] = 8'h30;
DFS[16'h2C39] = 8'h08;
DFS[16'h2C3A] = 8'hF0;
DFS[16'h2C3B] = 8'h03;
DFS[16'h2C3C] = 8'h4C;
DFS[16'h2C3D] = 8'h72;
DFS[16'h2C3E] = 8'hAA;
DFS[16'h2C3F] = 8'h4C;
DFS[16'h2C40] = 8'h78;
DFS[16'h2C41] = 8'hAA;
DFS[16'h2C42] = 8'hA8;
DFS[16'h2C43] = 8'hA9;
DFS[16'h2C44] = 8'hFF;
DFS[16'h2C45] = 8'h9D;
DFS[16'h2C46] = 8'h10;
DFS[16'h2C47] = 8'h0D;
DFS[16'h2C48] = 8'hC8;
DFS[16'h2C49] = 8'hD0;
DFS[16'h2C4A] = 8'h1A;
DFS[16'h2C4B] = 8'h20;
DFS[16'h2C4C] = 8'h00;
DFS[16'h2C4D] = 8'hA0;
DFS[16'h2C4E] = 8'hC7;
DFS[16'h2C4F] = 8'h44;
DFS[16'h2C50] = 8'h69;
DFS[16'h2C51] = 8'h73;
DFS[16'h2C52] = 8'h6B;
DFS[16'h2C53] = 8'h20;
DFS[16'h2C54] = 8'h6E;
DFS[16'h2C55] = 8'h75;
DFS[16'h2C56] = 8'h6D;
DFS[16'h2C57] = 8'h62;
DFS[16'h2C58] = 8'h65;
DFS[16'h2C59] = 8'h72;
DFS[16'h2C5A] = 8'h20;
DFS[16'h2C5B] = 8'h6E;
DFS[16'h2C5C] = 8'h6F;
DFS[16'h2C5D] = 8'h74;
DFS[16'h2C5E] = 8'h20;
DFS[16'h2C5F] = 8'h76;
DFS[16'h2C60] = 8'h61;
DFS[16'h2C61] = 8'h6C;
DFS[16'h2C62] = 8'h69;
DFS[16'h2C63] = 8'h64;
DFS[16'h2C64] = 8'h00;
DFS[16'h2C65] = 8'h20;
DFS[16'h2C66] = 8'h00;
DFS[16'h2C67] = 8'hA0;
DFS[16'h2C68] = 8'hC7;
DFS[16'h2C69] = 8'h44;
DFS[16'h2C6A] = 8'h69;
DFS[16'h2C6B] = 8'h73;
DFS[16'h2C6C] = 8'h6B;
DFS[16'h2C6D] = 8'h20;
DFS[16'h2C6E] = 8'h6E;
DFS[16'h2C6F] = 8'h6F;
DFS[16'h2C70] = 8'h74;
DFS[16'h2C71] = 8'h20;
DFS[16'h2C72] = 8'h66;
DFS[16'h2C73] = 8'h6F;
DFS[16'h2C74] = 8'h72;
DFS[16'h2C75] = 8'h6D;
DFS[16'h2C76] = 8'h61;
DFS[16'h2C77] = 8'h74;
DFS[16'h2C78] = 8'h74;
DFS[16'h2C79] = 8'h65;
DFS[16'h2C7A] = 8'h64;
DFS[16'h2C7B] = 8'h00;
DFS[16'h2C7C] = 8'h29;
DFS[16'h2C7D] = 8'h7E;
DFS[16'h2C7E] = 8'h48;
DFS[16'h2C7F] = 8'h20;
DFS[16'h2C80] = 8'h17;
DFS[16'h2C81] = 8'hA8;
DFS[16'h2C82] = 8'h18;
DFS[16'h2C83] = 8'h68;
DFS[16'h2C84] = 8'h6D;
DFS[16'h2C85] = 8'h06;
DFS[16'h2C86] = 8'h0D;
DFS[16'h2C87] = 8'h85;
DFS[16'h2C88] = 8'hA2;
DFS[16'h2C89] = 8'hAD;
DFS[16'h2C8A] = 8'h07;
DFS[16'h2C8B] = 8'h0D;
DFS[16'h2C8C] = 8'h69;
DFS[16'h2C8D] = 8'h00;
DFS[16'h2C8E] = 8'h85;
DFS[16'h2C8F] = 8'hA3;
DFS[16'h2C90] = 8'hAD;
DFS[16'h2C91] = 8'h08;
DFS[16'h2C92] = 8'h0D;
DFS[16'h2C93] = 8'h69;
DFS[16'h2C94] = 8'h00;
DFS[16'h2C95] = 8'h85;
DFS[16'h2C96] = 8'hA4;
DFS[16'h2C97] = 8'h60;
DFS[16'h2C98] = 8'h29;
DFS[16'h2C99] = 8'hFE;
DFS[16'h2C9A] = 8'h09;
DFS[16'h2C9B] = 8'h80;
DFS[16'h2C9C] = 8'hCD;
DFS[16'h2C9D] = 8'h82;
DFS[16'h2C9E] = 8'h10;
DFS[16'h2C9F] = 8'hF0;
DFS[16'h2CA0] = 8'hF6;
DFS[16'h2CA1] = 8'h8D;
DFS[16'h2CA2] = 8'h82;
DFS[16'h2CA3] = 8'h10;
DFS[16'h2CA4] = 8'h48;
DFS[16'h2CA5] = 8'h20;
DFS[16'h2CA6] = 8'hEC;
DFS[16'h2CA7] = 8'hA4;
DFS[16'h2CA8] = 8'h68;
DFS[16'h2CA9] = 8'h20;
DFS[16'h2CAA] = 8'h7C;
DFS[16'h2CAB] = 8'hAC;
DFS[16'h2CAC] = 8'h4C;
DFS[16'h2CAD] = 8'h0F;
DFS[16'h2CAE] = 8'hA6;
DFS[16'h2CAF] = 8'h8D;
DFS[16'h2CB0] = 8'h82;
DFS[16'h2CB1] = 8'h10;
DFS[16'h2CB2] = 8'h20;
DFS[16'h2CB3] = 8'h7C;
DFS[16'h2CB4] = 8'hAC;
DFS[16'h2CB5] = 8'h4C;
DFS[16'h2CB6] = 8'h0F;
DFS[16'h2CB7] = 8'hA6;
DFS[16'h2CB8] = 8'h20;
DFS[16'h2CB9] = 8'hEC;
DFS[16'h2CBA] = 8'hA4;
DFS[16'h2CBB] = 8'hAD;
DFS[16'h2CBC] = 8'h82;
DFS[16'h2CBD] = 8'h10;
DFS[16'h2CBE] = 8'h20;
DFS[16'h2CBF] = 8'h7C;
DFS[16'h2CC0] = 8'hAC;
DFS[16'h2CC1] = 8'h4C;
DFS[16'h2CC2] = 8'h28;
DFS[16'h2CC3] = 8'hA6;
DFS[16'h2CC4] = 8'hAD;
DFS[16'h2CC5] = 8'h82;
DFS[16'h2CC6] = 8'h10;
DFS[16'h2CC7] = 8'h20;
DFS[16'h2CC8] = 8'h7C;
DFS[16'h2CC9] = 8'hAC;
DFS[16'h2CCA] = 8'h4C;
DFS[16'h2CCB] = 8'h28;
DFS[16'h2CCC] = 8'hA6;
DFS[16'h2CCD] = 8'h20;
DFS[16'h2CCE] = 8'hB8;
DFS[16'h2CCF] = 8'hAC;
DFS[16'h2CD0] = 8'hA2;
DFS[16'h2CD1] = 8'h03;
DFS[16'h2CD2] = 8'h20;
DFS[16'h2CD3] = 8'hD9;
DFS[16'h2CD4] = 8'hAC;
DFS[16'h2CD5] = 8'hCA;
DFS[16'h2CD6] = 8'h10;
DFS[16'h2CD7] = 8'hFA;
DFS[16'h2CD8] = 8'h60;
DFS[16'h2CD9] = 8'hBD;
DFS[16'h2CDA] = 8'h10;
DFS[16'h2CDB] = 8'h0D;
DFS[16'h2CDC] = 8'h30;
DFS[16'h2CDD] = 8'h2B;
DFS[16'h2CDE] = 8'h49;
DFS[16'h2CDF] = 8'hFF;
DFS[16'h2CE0] = 8'hDD;
DFS[16'h2CE1] = 8'h18;
DFS[16'h2CE2] = 8'h0D;
DFS[16'h2CE3] = 8'hD0;
DFS[16'h2CE4] = 8'h18;
DFS[16'h2CE5] = 8'hBD;
DFS[16'h2CE6] = 8'h0C;
DFS[16'h2CE7] = 8'h0D;
DFS[16'h2CE8] = 8'h49;
DFS[16'h2CE9] = 8'hFF;
DFS[16'h2CEA] = 8'hDD;
DFS[16'h2CEB] = 8'h14;
DFS[16'h2CEC] = 8'h0D;
DFS[16'h2CED] = 8'hD0;
DFS[16'h2CEE] = 8'h0E;
DFS[16'h2CEF] = 8'hBD;
DFS[16'h2CF0] = 8'h10;
DFS[16'h2CF1] = 8'h0D;
DFS[16'h2CF2] = 8'h6A;
DFS[16'h2CF3] = 8'hBD;
DFS[16'h2CF4] = 8'h0C;
DFS[16'h2CF5] = 8'h0D;
DFS[16'h2CF6] = 8'h20;
DFS[16'h2CF7] = 8'hCD;
DFS[16'h2CF8] = 8'hAB;
DFS[16'h2CF9] = 8'hF0;
DFS[16'h2CFA] = 8'h0B;
DFS[16'h2CFB] = 8'h10;
DFS[16'h2CFC] = 8'h07;
DFS[16'h2CFD] = 8'hA9;
DFS[16'h2CFE] = 8'hFF;
DFS[16'h2CFF] = 8'h9D;
DFS[16'h2D00] = 8'h10;
DFS[16'h2D01] = 8'h0D;
DFS[16'h2D02] = 8'hD0;
DFS[16'h2D03] = 8'h02;
DFS[16'h2D04] = 8'hA9;
DFS[16'h2D05] = 8'h54;
DFS[16'h2D06] = 8'h9D;
DFS[16'h2D07] = 8'h1C;
DFS[16'h2D08] = 8'h0D;
DFS[16'h2D09] = 8'h60;
DFS[16'h2D0A] = 8'hA9;
DFS[16'h2D0B] = 8'hFF;
DFS[16'h2D0C] = 8'hA2;
DFS[16'h2D0D] = 8'h1F;
DFS[16'h2D0E] = 8'h9D;
DFS[16'h2D0F] = 8'h20;
DFS[16'h2D10] = 8'h0D;
DFS[16'h2D11] = 8'hCA;
DFS[16'h2D12] = 8'hD0;
DFS[16'h2D13] = 8'hFA;
DFS[16'h2D14] = 8'h8E;
DFS[16'h2D15] = 8'h04;
DFS[16'h2D16] = 8'h0D;
DFS[16'h2D17] = 8'hA9;
DFS[16'h2D18] = 8'h00;
DFS[16'h2D19] = 8'h8D;
DFS[16'h2D1A] = 8'h02;
DFS[16'h2D1B] = 8'h0D;
DFS[16'h2D1C] = 8'h8D;
DFS[16'h2D1D] = 8'h05;
DFS[16'h2D1E] = 8'h0D;
DFS[16'h2D1F] = 8'h8D;
DFS[16'h2D20] = 8'h20;
DFS[16'h2D21] = 8'h0D;
DFS[16'h2D22] = 8'hA9;
DFS[16'h2D23] = 8'h80;
DFS[16'h2D24] = 8'h20;
DFS[16'h2D25] = 8'hA1;
DFS[16'h2D26] = 8'hAC;
DFS[16'h2D27] = 8'hA2;
DFS[16'h2D28] = 8'h00;
DFS[16'h2D29] = 8'hAD;
DFS[16'h2D2A] = 8'h52;
DFS[16'h2D2B] = 8'h0D;
DFS[16'h2D2C] = 8'hC9;
DFS[16'h2D2D] = 8'h42;
DFS[16'h2D2E] = 8'hF0;
DFS[16'h2D2F] = 8'h16;
DFS[16'h2D30] = 8'hBD;
DFS[16'h2D31] = 8'h10;
DFS[16'h2D32] = 8'h0D;
DFS[16'h2D33] = 8'h30;
DFS[16'h2D34] = 8'h43;
DFS[16'h2D35] = 8'h49;
DFS[16'h2D36] = 8'hFF;
DFS[16'h2D37] = 8'hDD;
DFS[16'h2D38] = 8'h18;
DFS[16'h2D39] = 8'h0D;
DFS[16'h2D3A] = 8'hD0;
DFS[16'h2D3B] = 8'h0A;
DFS[16'h2D3C] = 8'hBD;
DFS[16'h2D3D] = 8'h0C;
DFS[16'h2D3E] = 8'h0D;
DFS[16'h2D3F] = 8'h49;
DFS[16'h2D40] = 8'hFF;
DFS[16'h2D41] = 8'hDD;
DFS[16'h2D42] = 8'h14;
DFS[16'h2D43] = 8'h0D;
DFS[16'h2D44] = 8'hF0;
DFS[16'h2D45] = 8'h16;
DFS[16'h2D46] = 8'hBD;
DFS[16'h2D47] = 8'h00;
DFS[16'h2D48] = 8'h0E;
DFS[16'h2D49] = 8'h9D;
DFS[16'h2D4A] = 8'h0C;
DFS[16'h2D4B] = 8'h0D;
DFS[16'h2D4C] = 8'h49;
DFS[16'h2D4D] = 8'hFF;
DFS[16'h2D4E] = 8'h9D;
DFS[16'h2D4F] = 8'h14;
DFS[16'h2D50] = 8'h0D;
DFS[16'h2D51] = 8'hBD;
DFS[16'h2D52] = 8'h04;
DFS[16'h2D53] = 8'h0E;
DFS[16'h2D54] = 8'h9D;
DFS[16'h2D55] = 8'h10;
DFS[16'h2D56] = 8'h0D;
DFS[16'h2D57] = 8'h49;
DFS[16'h2D58] = 8'hFF;
DFS[16'h2D59] = 8'h9D;
DFS[16'h2D5A] = 8'h18;
DFS[16'h2D5B] = 8'h0D;
DFS[16'h2D5C] = 8'h8A;
DFS[16'h2D5D] = 8'hF0;
DFS[16'h2D5E] = 8'h1E;
DFS[16'h2D5F] = 8'hA8;
DFS[16'h2D60] = 8'h88;
DFS[16'h2D61] = 8'hBD;
DFS[16'h2D62] = 8'h10;
DFS[16'h2D63] = 8'h0D;
DFS[16'h2D64] = 8'h30;
DFS[16'h2D65] = 8'h17;
DFS[16'h2D66] = 8'hD9;
DFS[16'h2D67] = 8'h10;
DFS[16'h2D68] = 8'h0D;
DFS[16'h2D69] = 8'hD0;
DFS[16'h2D6A] = 8'h08;
DFS[16'h2D6B] = 8'hBD;
DFS[16'h2D6C] = 8'h0C;
DFS[16'h2D6D] = 8'h0D;
DFS[16'h2D6E] = 8'hD9;
DFS[16'h2D6F] = 8'h0C;
DFS[16'h2D70] = 8'h0D;
DFS[16'h2D71] = 8'hF0;
DFS[16'h2D72] = 8'h05;
DFS[16'h2D73] = 8'h88;
DFS[16'h2D74] = 8'h10;
DFS[16'h2D75] = 8'hEB;
DFS[16'h2D76] = 8'h30;
DFS[16'h2D77] = 8'h05;
DFS[16'h2D78] = 8'hA9;
DFS[16'h2D79] = 8'hFF;
DFS[16'h2D7A] = 8'h9D;
DFS[16'h2D7B] = 8'h10;
DFS[16'h2D7C] = 8'h0D;
DFS[16'h2D7D] = 8'hE8;
DFS[16'h2D7E] = 8'hE0;
DFS[16'h2D7F] = 8'h04;
DFS[16'h2D80] = 8'hD0;
DFS[16'h2D81] = 8'hA7;
DFS[16'h2D82] = 8'h4C;
DFS[16'h2D83] = 8'hD0;
DFS[16'h2D84] = 8'hAC;
DFS[16'h2D85] = 8'h08;
DFS[16'h2D86] = 8'h48;
DFS[16'h2D87] = 8'h8D;
DFS[16'h2D88] = 8'h53;
DFS[16'h2D89] = 8'h0D;
DFS[16'h2D8A] = 8'hA9;
DFS[16'h2D8B] = 8'h00;
DFS[16'h2D8C] = 8'h2A;
DFS[16'h2D8D] = 8'h8D;
DFS[16'h2D8E] = 8'h54;
DFS[16'h2D8F] = 8'h0D;
DFS[16'h2D90] = 8'h68;
DFS[16'h2D91] = 8'h28;
DFS[16'h2D92] = 8'h08;
DFS[16'h2D93] = 8'h48;
DFS[16'h2D94] = 8'h20;
DFS[16'h2D95] = 8'hCD;
DFS[16'h2D96] = 8'hA9;
DFS[16'h2D97] = 8'h8E;
DFS[16'h2D98] = 8'h55;
DFS[16'h2D99] = 8'h0D;
DFS[16'h2D9A] = 8'h8D;
DFS[16'h2D9B] = 8'h56;
DFS[16'h2D9C] = 8'h0D;
DFS[16'h2D9D] = 8'h68;
DFS[16'h2D9E] = 8'h28;
DFS[16'h2D9F] = 8'h20;
DFS[16'h2DA0] = 8'hB9;
DFS[16'h2DA1] = 8'hAB;
DFS[16'h2DA2] = 8'h29;
DFS[16'h2DA3] = 8'hF0;
DFS[16'h2DA4] = 8'h85;
DFS[16'h2DA5] = 8'hF2;
DFS[16'h2DA6] = 8'h98;
DFS[16'h2DA7] = 8'h29;
DFS[16'h2DA8] = 8'h01;
DFS[16'h2DA9] = 8'h09;
DFS[16'h2DAA] = 8'h0E;
DFS[16'h2DAB] = 8'h85;
DFS[16'h2DAC] = 8'hF3;
DFS[16'h2DAD] = 8'h98;
DFS[16'h2DAE] = 8'h29;
DFS[16'h2DAF] = 8'hFE;
DFS[16'h2DB0] = 8'h09;
DFS[16'h2DB1] = 8'h80;
DFS[16'h2DB2] = 8'h8D;
DFS[16'h2DB3] = 8'h52;
DFS[16'h2DB4] = 8'h0D;
DFS[16'h2DB5] = 8'h20;
DFS[16'h2DB6] = 8'h9C;
DFS[16'h2DB7] = 8'hAC;
DFS[16'h2DB8] = 8'h4C;
DFS[16'h2DB9] = 8'h19;
DFS[16'h2DBA] = 8'hAE;
DFS[16'h2DBB] = 8'hA9;
DFS[16'h2DBC] = 8'h00;
DFS[16'h2DBD] = 8'h8D;
DFS[16'h2DBE] = 8'h55;
DFS[16'h2DBF] = 8'h0D;
DFS[16'h2DC0] = 8'h8D;
DFS[16'h2DC1] = 8'h56;
DFS[16'h2DC2] = 8'h0D;
DFS[16'h2DC3] = 8'h8D;
DFS[16'h2DC4] = 8'h53;
DFS[16'h2DC5] = 8'h0D;
DFS[16'h2DC6] = 8'h8D;
DFS[16'h2DC7] = 8'h54;
DFS[16'h2DC8] = 8'h0D;
DFS[16'h2DC9] = 8'hA9;
DFS[16'h2DCA] = 8'h10;
DFS[16'h2DCB] = 8'h85;
DFS[16'h2DCC] = 8'hF2;
DFS[16'h2DCD] = 8'hA9;
DFS[16'h2DCE] = 8'h0E;
DFS[16'h2DCF] = 8'h85;
DFS[16'h2DD0] = 8'hF3;
DFS[16'h2DD1] = 8'hA9;
DFS[16'h2DD2] = 8'h80;
DFS[16'h2DD3] = 8'h8D;
DFS[16'h2DD4] = 8'h52;
DFS[16'h2DD5] = 8'h0D;
DFS[16'h2DD6] = 8'h20;
DFS[16'h2DD7] = 8'h9C;
DFS[16'h2DD8] = 8'hAC;
DFS[16'h2DD9] = 8'h4C;
DFS[16'h2DDA] = 8'h19;
DFS[16'h2DDB] = 8'hAE;
DFS[16'h2DDC] = 8'hC9;
DFS[16'h2DDD] = 8'hFF;
DFS[16'h2DDE] = 8'hF0;
DFS[16'h2DDF] = 8'h41;
DFS[16'h2DE0] = 8'h18;
DFS[16'h2DE1] = 8'hA5;
DFS[16'h2DE2] = 8'hF2;
DFS[16'h2DE3] = 8'h69;
DFS[16'h2DE4] = 8'h10;
DFS[16'h2DE5] = 8'h85;
DFS[16'h2DE6] = 8'hF2;
DFS[16'h2DE7] = 8'hD0;
DFS[16'h2DE8] = 8'h18;
DFS[16'h2DE9] = 8'hA5;
DFS[16'h2DEA] = 8'hF3;
DFS[16'h2DEB] = 8'h49;
DFS[16'h2DEC] = 8'h01;
DFS[16'h2DED] = 8'h85;
DFS[16'h2DEE] = 8'hF3;
DFS[16'h2DEF] = 8'h6A;
DFS[16'h2DF0] = 8'hB0;
DFS[16'h2DF1] = 8'h0F;
DFS[16'h2DF2] = 8'hAD;
DFS[16'h2DF3] = 8'h52;
DFS[16'h2DF4] = 8'h0D;
DFS[16'h2DF5] = 8'h69;
DFS[16'h2DF6] = 8'h02;
DFS[16'h2DF7] = 8'hC9;
DFS[16'h2DF8] = 8'hA0;
DFS[16'h2DF9] = 8'hF0;
DFS[16'h2DFA] = 8'h26;
DFS[16'h2DFB] = 8'h8D;
DFS[16'h2DFC] = 8'h52;
DFS[16'h2DFD] = 8'h0D;
DFS[16'h2DFE] = 8'h20;
DFS[16'h2DFF] = 8'h9C;
DFS[16'h2E00] = 8'hAC;
DFS[16'h2E01] = 8'hEE;
DFS[16'h2E02] = 8'h53;
DFS[16'h2E03] = 8'h0D;
DFS[16'h2E04] = 8'hD0;
DFS[16'h2E05] = 8'h03;
DFS[16'h2E06] = 8'hEE;
DFS[16'h2E07] = 8'h54;
DFS[16'h2E08] = 8'h0D;
DFS[16'h2E09] = 8'hF8;
DFS[16'h2E0A] = 8'h18;
DFS[16'h2E0B] = 8'hAD;
DFS[16'h2E0C] = 8'h55;
DFS[16'h2E0D] = 8'h0D;
DFS[16'h2E0E] = 8'h69;
DFS[16'h2E0F] = 8'h01;
DFS[16'h2E10] = 8'h8D;
DFS[16'h2E11] = 8'h55;
DFS[16'h2E12] = 8'h0D;
DFS[16'h2E13] = 8'h90;
DFS[16'h2E14] = 8'h03;
DFS[16'h2E15] = 8'hEE;
DFS[16'h2E16] = 8'h56;
DFS[16'h2E17] = 8'h0D;
DFS[16'h2E18] = 8'hD8;
DFS[16'h2E19] = 8'hA0;
DFS[16'h2E1A] = 8'h0F;
DFS[16'h2E1B] = 8'hB1;
DFS[16'h2E1C] = 8'hF2;
DFS[16'h2E1D] = 8'h30;
DFS[16'h2E1E] = 8'hBD;
DFS[16'h2E1F] = 8'h18;
DFS[16'h2E20] = 8'h60;
DFS[16'h2E21] = 8'hA9;
DFS[16'h2E22] = 8'hFF;
DFS[16'h2E23] = 8'h8D;
DFS[16'h2E24] = 8'h54;
DFS[16'h2E25] = 8'h0D;
DFS[16'h2E26] = 8'h38;
DFS[16'h2E27] = 8'h60;
DFS[16'h2E28] = 8'h20;
DFS[16'h2E29] = 8'hEC;
DFS[16'h2E2A] = 8'hA4;
DFS[16'h2E2B] = 8'hA9;
DFS[16'h2E2C] = 8'h80;
DFS[16'h2E2D] = 8'h8D;
DFS[16'h2E2E] = 8'h52;
DFS[16'h2E2F] = 8'h0D;
DFS[16'h2E30] = 8'h20;
DFS[16'h2E31] = 8'hAF;
DFS[16'h2E32] = 8'hAC;
DFS[16'h2E33] = 8'hA9;
DFS[16'h2E34] = 8'h10;
DFS[16'h2E35] = 8'h85;
DFS[16'h2E36] = 8'hF2;
DFS[16'h2E37] = 8'hA9;
DFS[16'h2E38] = 8'h0E;
DFS[16'h2E39] = 8'h85;
DFS[16'h2E3A] = 8'hF3;
DFS[16'h2E3B] = 8'h20;
DFS[16'h2E3C] = 8'h17;
DFS[16'h2E3D] = 8'hA8;
DFS[16'h2E3E] = 8'h18;
DFS[16'h2E3F] = 8'hAD;
DFS[16'h2E40] = 8'h06;
DFS[16'h2E41] = 8'h0D;
DFS[16'h2E42] = 8'h69;
DFS[16'h2E43] = 8'h20;
DFS[16'h2E44] = 8'h85;
DFS[16'h2E45] = 8'hA2;
DFS[16'h2E46] = 8'hAD;
DFS[16'h2E47] = 8'h07;
DFS[16'h2E48] = 8'h0D;
DFS[16'h2E49] = 8'h69;
DFS[16'h2E4A] = 8'h00;
DFS[16'h2E4B] = 8'h85;
DFS[16'h2E4C] = 8'hA3;
DFS[16'h2E4D] = 8'hAD;
DFS[16'h2E4E] = 8'h08;
DFS[16'h2E4F] = 8'h0D;
DFS[16'h2E50] = 8'h69;
DFS[16'h2E51] = 8'h00;
DFS[16'h2E52] = 8'h85;
DFS[16'h2E53] = 8'hA4;
DFS[16'h2E54] = 8'h20;
DFS[16'h2E55] = 8'h9B;
DFS[16'h2E56] = 8'hA7;
DFS[16'h2E57] = 8'hA0;
DFS[16'h2E58] = 8'h0F;
DFS[16'h2E59] = 8'hB1;
DFS[16'h2E5A] = 8'hF2;
DFS[16'h2E5B] = 8'hC9;
DFS[16'h2E5C] = 8'hFF;
DFS[16'h2E5D] = 8'hF0;
DFS[16'h2E5E] = 8'h39;
DFS[16'h2E5F] = 8'h20;
DFS[16'h2E60] = 8'hB2;
DFS[16'h2E61] = 8'hA7;
DFS[16'h2E62] = 8'hA0;
DFS[16'h2E63] = 8'h0B;
DFS[16'h2E64] = 8'hB9;
DFS[16'h2E65] = 8'h5F;
DFS[16'h2E66] = 8'h0D;
DFS[16'h2E67] = 8'h91;
DFS[16'h2E68] = 8'hF2;
DFS[16'h2E69] = 8'h88;
DFS[16'h2E6A] = 8'h10;
DFS[16'h2E6B] = 8'hF8;
DFS[16'h2E6C] = 8'h18;
DFS[16'h2E6D] = 8'hA5;
DFS[16'h2E6E] = 8'hF2;
DFS[16'h2E6F] = 8'h69;
DFS[16'h2E70] = 8'h10;
DFS[16'h2E71] = 8'h85;
DFS[16'h2E72] = 8'hF2;
DFS[16'h2E73] = 8'hD0;
DFS[16'h2E74] = 8'hE2;
DFS[16'h2E75] = 8'hA5;
DFS[16'h2E76] = 8'hF3;
DFS[16'h2E77] = 8'h49;
DFS[16'h2E78] = 8'h01;
DFS[16'h2E79] = 8'h85;
DFS[16'h2E7A] = 8'hF3;
DFS[16'h2E7B] = 8'h6A;
DFS[16'h2E7C] = 8'hB0;
DFS[16'h2E7D] = 8'hD9;
DFS[16'h2E7E] = 8'h20;
DFS[16'h2E7F] = 8'hC4;
DFS[16'h2E80] = 8'hAC;
DFS[16'h2E81] = 8'h18;
DFS[16'h2E82] = 8'hAD;
DFS[16'h2E83] = 8'h52;
DFS[16'h2E84] = 8'h0D;
DFS[16'h2E85] = 8'h69;
DFS[16'h2E86] = 8'h02;
DFS[16'h2E87] = 8'hC9;
DFS[16'h2E88] = 8'hA0;
DFS[16'h2E89] = 8'hF0;
DFS[16'h2E8A] = 8'h18;
DFS[16'h2E8B] = 8'h8D;
DFS[16'h2E8C] = 8'h52;
DFS[16'h2E8D] = 8'h0D;
DFS[16'h2E8E] = 8'h24;
DFS[16'h2E8F] = 8'hFF;
DFS[16'h2E90] = 8'h30;
DFS[16'h2E91] = 8'h12;
DFS[16'h2E92] = 8'h20;
DFS[16'h2E93] = 8'hAF;
DFS[16'h2E94] = 8'hAC;
DFS[16'h2E95] = 8'h4C;
DFS[16'h2E96] = 8'h57;
DFS[16'h2E97] = 8'hAE;
DFS[16'h2E98] = 8'hA5;
DFS[16'h2E99] = 8'hF2;
DFS[16'h2E9A] = 8'hD0;
DFS[16'h2E9B] = 8'h04;
DFS[16'h2E9C] = 8'h66;
DFS[16'h2E9D] = 8'hF3;
DFS[16'h2E9E] = 8'h90;
DFS[16'h2E9F] = 8'h03;
DFS[16'h2EA0] = 8'h20;
DFS[16'h2EA1] = 8'hC4;
DFS[16'h2EA2] = 8'hAC;
DFS[16'h2EA3] = 8'h60;
DFS[16'h2EA4] = 8'h4C;
DFS[16'h2EA5] = 8'h82;
DFS[16'h2EA6] = 8'hA0;
DFS[16'h2EA7] = 8'hA2;
DFS[16'h2EA8] = 8'h0B;
DFS[16'h2EA9] = 8'hA9;
DFS[16'h2EAA] = 8'h00;
DFS[16'h2EAB] = 8'h20;
DFS[16'h2EAC] = 8'hC6;
DFS[16'h2EAD] = 8'h88;
DFS[16'h2EAE] = 8'h9D;
DFS[16'h2EAF] = 8'h5F;
DFS[16'h2EB0] = 8'h0D;
DFS[16'h2EB1] = 8'hCA;
DFS[16'h2EB2] = 8'h10;
DFS[16'h2EB3] = 8'hF7;
DFS[16'h2EB4] = 8'hE8;
DFS[16'h2EB5] = 8'h20;
DFS[16'h2EB6] = 8'hC5;
DFS[16'h2EB7] = 8'hFF;
DFS[16'h2EB8] = 8'hB0;
DFS[16'h2EB9] = 8'h0A;
DFS[16'h2EBA] = 8'h20;
DFS[16'h2EBB] = 8'hC6;
DFS[16'h2EBC] = 8'h88;
DFS[16'h2EBD] = 8'h9D;
DFS[16'h2EBE] = 8'h5F;
DFS[16'h2EBF] = 8'h0D;
DFS[16'h2EC0] = 8'hE0;
DFS[16'h2EC1] = 8'h0B;
DFS[16'h2EC2] = 8'h90;
DFS[16'h2EC3] = 8'hF0;
DFS[16'h2EC4] = 8'h20;
DFS[16'h2EC5] = 8'hB4;
DFS[16'h2EC6] = 8'h8A;
DFS[16'h2EC7] = 8'hAE;
DFS[16'h2EC8] = 8'h82;
DFS[16'h2EC9] = 8'h10;
DFS[16'h2ECA] = 8'hBD;
DFS[16'h2ECB] = 8'h10;
DFS[16'h2ECC] = 8'h0D;
DFS[16'h2ECD] = 8'h6A;
DFS[16'h2ECE] = 8'hBD;
DFS[16'h2ECF] = 8'h0C;
DFS[16'h2ED0] = 8'h0D;
DFS[16'h2ED1] = 8'h20;
DFS[16'h2ED2] = 8'hB9;
DFS[16'h2ED3] = 8'hAB;
DFS[16'h2ED4] = 8'h29;
DFS[16'h2ED5] = 8'hF0;
DFS[16'h2ED6] = 8'h48;
DFS[16'h2ED7] = 8'h98;
DFS[16'h2ED8] = 8'h48;
DFS[16'h2ED9] = 8'h29;
DFS[16'h2EDA] = 8'hFE;
DFS[16'h2EDB] = 8'h09;
DFS[16'h2EDC] = 8'h80;
DFS[16'h2EDD] = 8'h20;
DFS[16'h2EDE] = 8'hA1;
DFS[16'h2EDF] = 8'hAC;
DFS[16'h2EE0] = 8'h68;
DFS[16'h2EE1] = 8'h18;
DFS[16'h2EE2] = 8'h29;
DFS[16'h2EE3] = 8'h01;
DFS[16'h2EE4] = 8'h69;
DFS[16'h2EE5] = 8'h0E;
DFS[16'h2EE6] = 8'h85;
DFS[16'h2EE7] = 8'hF3;
DFS[16'h2EE8] = 8'h68;
DFS[16'h2EE9] = 8'h85;
DFS[16'h2EEA] = 8'hF2;
DFS[16'h2EEB] = 8'hA0;
DFS[16'h2EEC] = 8'h0B;
DFS[16'h2EED] = 8'hB9;
DFS[16'h2EEE] = 8'h5F;
DFS[16'h2EEF] = 8'h0D;
DFS[16'h2EF0] = 8'h91;
DFS[16'h2EF1] = 8'hF2;
DFS[16'h2EF2] = 8'h88;
DFS[16'h2EF3] = 8'h10;
DFS[16'h2EF4] = 8'hF8;
DFS[16'h2EF5] = 8'h4C;
DFS[16'h2EF6] = 8'hB8;
DFS[16'h2EF7] = 8'hAC;
DFS[16'h2EF8] = 8'h44;
DFS[16'h2EF9] = 8'h49;
DFS[16'h2EFA] = 8'h4E;
DFS[16'h2EFB] = 8'hB3;
DFS[16'h2EFC] = 8'hC0;
DFS[16'h2EFD] = 8'h12;
DFS[16'h2EFE] = 8'h44;
DFS[16'h2EFF] = 8'h42;
DFS[16'h2F00] = 8'h4F;
DFS[16'h2F01] = 8'h4F;
DFS[16'h2F02] = 8'h54;
DFS[16'h2F03] = 8'hB3;
DFS[16'h2F04] = 8'hB5;
DFS[16'h2F05] = 8'h02;
DFS[16'h2F06] = 8'h44;
DFS[16'h2F07] = 8'h43;
DFS[16'h2F08] = 8'h41;
DFS[16'h2F09] = 8'h54;
DFS[16'h2F0A] = 8'hB3;
DFS[16'h2F0B] = 8'hC6;
DFS[16'h2F0C] = 8'h04;
DFS[16'h2F0D] = 8'h44;
DFS[16'h2F0E] = 8'h44;
DFS[16'h2F0F] = 8'h49;
DFS[16'h2F10] = 8'h53;
DFS[16'h2F11] = 8'h4B;
DFS[16'h2F12] = 8'h53;
DFS[16'h2F13] = 8'hB5;
DFS[16'h2F14] = 8'h76;
DFS[16'h2F15] = 8'h01;
DFS[16'h2F16] = 8'h44;
DFS[16'h2F17] = 8'h4C;
DFS[16'h2F18] = 8'h4F;
DFS[16'h2F19] = 8'h43;
DFS[16'h2F1A] = 8'h4B;
DFS[16'h2F1B] = 8'hB5;
DFS[16'h2F1C] = 8'hBC;
DFS[16'h2F1D] = 8'h02;
DFS[16'h2F1E] = 8'h44;
DFS[16'h2F1F] = 8'h55;
DFS[16'h2F20] = 8'h4E;
DFS[16'h2F21] = 8'h4C;
DFS[16'h2F22] = 8'h4F;
DFS[16'h2F23] = 8'h43;
DFS[16'h2F24] = 8'h4B;
DFS[16'h2F25] = 8'hB5;
DFS[16'h2F26] = 8'hC0;
DFS[16'h2F27] = 8'h02;
DFS[16'h2F28] = 8'h44;
DFS[16'h2F29] = 8'h46;
DFS[16'h2F2A] = 8'h52;
DFS[16'h2F2B] = 8'h45;
DFS[16'h2F2C] = 8'h45;
DFS[16'h2F2D] = 8'hB4;
DFS[16'h2F2E] = 8'hB0;
DFS[16'h2F2F] = 8'h00;
DFS[16'h2F30] = 8'h44;
DFS[16'h2F31] = 8'h4B;
DFS[16'h2F32] = 8'h49;
DFS[16'h2F33] = 8'h4C;
DFS[16'h2F34] = 8'h4C;
DFS[16'h2F35] = 8'hB5;
DFS[16'h2F36] = 8'hE3;
DFS[16'h2F37] = 8'h03;
DFS[16'h2F38] = 8'h44;
DFS[16'h2F39] = 8'h52;
DFS[16'h2F3A] = 8'h45;
DFS[16'h2F3B] = 8'h53;
DFS[16'h2F3C] = 8'h54;
DFS[16'h2F3D] = 8'h4F;
DFS[16'h2F3E] = 8'h52;
DFS[16'h2F3F] = 8'h45;
DFS[16'h2F40] = 8'hB6;
DFS[16'h2F41] = 8'h26;
DFS[16'h2F42] = 8'h03;
DFS[16'h2F43] = 8'h44;
DFS[16'h2F44] = 8'h4E;
DFS[16'h2F45] = 8'h45;
DFS[16'h2F46] = 8'h57;
DFS[16'h2F47] = 8'hB6;
DFS[16'h2F48] = 8'h7B;
DFS[16'h2F49] = 8'h01;
DFS[16'h2F4A] = 8'h44;
DFS[16'h2F4B] = 8'h46;
DFS[16'h2F4C] = 8'h4F;
DFS[16'h2F4D] = 8'h52;
DFS[16'h2F4E] = 8'h4D;
DFS[16'h2F4F] = 8'hB6;
DFS[16'h2F50] = 8'h1E;
DFS[16'h2F51] = 8'h03;
DFS[16'h2F52] = 8'h44;
DFS[16'h2F53] = 8'h4F;
DFS[16'h2F54] = 8'h4E;
DFS[16'h2F55] = 8'h42;
DFS[16'h2F56] = 8'h4F;
DFS[16'h2F57] = 8'h4F;
DFS[16'h2F58] = 8'h54;
DFS[16'h2F59] = 8'hB7;
DFS[16'h2F5A] = 8'h49;
DFS[16'h2F5B] = 8'h52;
DFS[16'h2F5C] = 8'h44;
DFS[16'h2F5D] = 8'h52;
DFS[16'h2F5E] = 8'h45;
DFS[16'h2F5F] = 8'h43;
DFS[16'h2F60] = 8'h41;
DFS[16'h2F61] = 8'h54;
DFS[16'h2F62] = 8'hAE;
DFS[16'h2F63] = 8'h27;
DFS[16'h2F64] = 8'h00;
DFS[16'h2F65] = 8'h44;
DFS[16'h2F66] = 8'h52;
DFS[16'h2F67] = 8'h4F;
DFS[16'h2F68] = 8'h4D;
DFS[16'h2F69] = 8'hB7;
DFS[16'h2F6A] = 8'hB0;
DFS[16'h2F6B] = 8'h86;
DFS[16'h2F6C] = 8'h44;
DFS[16'h2F6D] = 8'h4D;
DFS[16'h2F6E] = 8'h4F;
DFS[16'h2F6F] = 8'h44;
DFS[16'h2F70] = 8'h45;
DFS[16'h2F71] = 8'hB7;
DFS[16'h2F72] = 8'h64;
DFS[16'h2F73] = 8'h07;
DFS[16'h2F74] = 8'h44;
DFS[16'h2F75] = 8'h53;
DFS[16'h2F76] = 8'h57;
DFS[16'h2F77] = 8'h41;
DFS[16'h2F78] = 8'h50;
DFS[16'h2F79] = 8'hB7;
DFS[16'h2F7A] = 8'h9A;
DFS[16'h2F7B] = 8'h00;
DFS[16'h2F7C] = 8'h44;
DFS[16'h2F7D] = 8'h41;
DFS[16'h2F7E] = 8'h42;
DFS[16'h2F7F] = 8'h4F;
DFS[16'h2F80] = 8'h55;
DFS[16'h2F81] = 8'h54;
DFS[16'h2F82] = 8'hAF;
DFS[16'h2F83] = 8'hFA;
DFS[16'h2F84] = 8'h00;
DFS[16'h2F85] = 8'h87;
DFS[16'h2F86] = 8'hD6;
DFS[16'h2F87] = 8'h00;
DFS[16'h2F88] = 8'h44;
DFS[16'h2F89] = 8'h55;
DFS[16'h2F8A] = 8'h54;
DFS[16'h2F8B] = 8'h49;
DFS[16'h2F8C] = 8'h4C;
DFS[16'h2F8D] = 8'h53;
DFS[16'h2F8E] = 8'hAF;
DFS[16'h2F8F] = 8'hCB;
DFS[16'h2F90] = 8'h00;
DFS[16'h2F91] = 8'hAF;
DFS[16'h2F92] = 8'hBD;
DFS[16'h2F93] = 8'h00;
DFS[16'h2F94] = 8'hA2;
DFS[16'h2F95] = 8'hA0;
DFS[16'h2F96] = 8'hB1;
DFS[16'h2F97] = 8'hF2;
DFS[16'h2F98] = 8'hC9;
DFS[16'h2F99] = 8'h0D;
DFS[16'h2F9A] = 8'hD0;
DFS[16'h2F9B] = 8'h16;
DFS[16'h2F9C] = 8'h98;
DFS[16'h2F9D] = 8'hE8;
DFS[16'h2F9E] = 8'hA0;
DFS[16'h2F9F] = 8'h02;
DFS[16'h2FA0] = 8'h20;
DFS[16'h2FA1] = 8'hCB;
DFS[16'h2FA2] = 8'h99;
DFS[16'h2FA3] = 8'h20;
DFS[16'h2FA4] = 8'hFF;
DFS[16'h2FA5] = 8'hB1;
DFS[16'h2FA6] = 8'h20;
DFS[16'h2FA7] = 8'h20;
DFS[16'h2FA8] = 8'h44;
DFS[16'h2FA9] = 8'h55;
DFS[16'h2FAA] = 8'h54;
DFS[16'h2FAB] = 8'h49;
DFS[16'h2FAC] = 8'h4C;
DFS[16'h2FAD] = 8'h53;
DFS[16'h2FAE] = 8'h00;
DFS[16'h2FAF] = 8'h4C;
DFS[16'h2FB0] = 8'hE7;
DFS[16'h2FB1] = 8'hFF;
DFS[16'h2FB2] = 8'h98;
DFS[16'h2FB3] = 8'h48;
DFS[16'h2FB4] = 8'h20;
DFS[16'h2FB5] = 8'h71;
DFS[16'h2FB6] = 8'h86;
DFS[16'h2FB7] = 8'h68;
DFS[16'h2FB8] = 8'hA8;
DFS[16'h2FB9] = 8'hA2;
DFS[16'h2FBA] = 8'h8D;
DFS[16'h2FBB] = 8'h4C;
DFS[16'h2FBC] = 8'h29;
DFS[16'h2FBD] = 8'hB0;
DFS[16'h2FBE] = 8'hC8;
DFS[16'h2FBF] = 8'hB1;
DFS[16'h2FC0] = 8'hF2;
DFS[16'h2FC1] = 8'hC9;
DFS[16'h2FC2] = 8'h0D;
DFS[16'h2FC3] = 8'hF0;
DFS[16'h2FC4] = 8'h06;
DFS[16'h2FC5] = 8'hC9;
DFS[16'h2FC6] = 8'h20;
DFS[16'h2FC7] = 8'hF0;
DFS[16'h2FC8] = 8'hF0;
DFS[16'h2FC9] = 8'hD0;
DFS[16'h2FCA] = 8'hF3;
DFS[16'h2FCB] = 8'h60;
DFS[16'h2FCC] = 8'h20;
DFS[16'h2FCD] = 8'hE7;
DFS[16'h2FCE] = 8'hFF;
DFS[16'h2FCF] = 8'h20;
DFS[16'h2FD0] = 8'hFF;
DFS[16'h2FD1] = 8'hB1;
DFS[16'h2FD2] = 8'h44;
DFS[16'h2FD3] = 8'h46;
DFS[16'h2FD4] = 8'h53;
DFS[16'h2FD5] = 8'h20;
DFS[16'h2FD6] = 8'h30;
DFS[16'h2FD7] = 8'h2E;
DFS[16'h2FD8] = 8'h39;
DFS[16'h2FD9] = 8'h30;
DFS[16'h2FDA] = 8'h00;
DFS[16'h2FDB] = 8'h20;
DFS[16'h2FDC] = 8'hE7;
DFS[16'h2FDD] = 8'hFF;
DFS[16'h2FDE] = 8'hA2;
DFS[16'h2FDF] = 8'h00;
DFS[16'h2FE0] = 8'hA9;
DFS[16'h2FE1] = 8'h0E;
DFS[16'h2FE2] = 8'h86;
DFS[16'h2FE3] = 8'hB5;
DFS[16'h2FE4] = 8'h85;
DFS[16'h2FE5] = 8'hBF;
DFS[16'h2FE6] = 8'hA2;
DFS[16'h2FE7] = 8'h00;
DFS[16'h2FE8] = 8'hA9;
DFS[16'h2FE9] = 8'h20;
DFS[16'h2FEA] = 8'h20;
DFS[16'h2FEB] = 8'hEE;
DFS[16'h2FEC] = 8'hFF;
DFS[16'h2FED] = 8'h20;
DFS[16'h2FEE] = 8'hEE;
DFS[16'h2FEF] = 8'hFF;
DFS[16'h2FF0] = 8'h20;
DFS[16'h2FF1] = 8'hC3;
DFS[16'h2FF2] = 8'hB2;
DFS[16'h2FF3] = 8'h20;
DFS[16'h2FF4] = 8'hE7;
DFS[16'h2FF5] = 8'hFF;
DFS[16'h2FF6] = 8'hC6;
DFS[16'h2FF7] = 8'hBF;
DFS[16'h2FF8] = 8'hD0;
DFS[16'h2FF9] = 8'hEE;
DFS[16'h2FFA] = 8'h60;
DFS[16'h2FFB] = 8'h20;
DFS[16'h2FFC] = 8'hFF;
DFS[16'h2FFD] = 8'hB1;
DFS[16'h2FFE] = 8'h44;
DFS[16'h2FFF] = 8'h55;
DFS[16'h3000] = 8'h54;
DFS[16'h3001] = 8'h49;
DFS[16'h3002] = 8'h4C;
DFS[16'h3003] = 8'h53;
DFS[16'h3004] = 8'h20;
DFS[16'h3005] = 8'h62;
DFS[16'h3006] = 8'h79;
DFS[16'h3007] = 8'h20;
DFS[16'h3008] = 8'h4D;
DFS[16'h3009] = 8'h61;
DFS[16'h300A] = 8'h72;
DFS[16'h300B] = 8'h74;
DFS[16'h300C] = 8'h69;
DFS[16'h300D] = 8'h6E;
DFS[16'h300E] = 8'h20;
DFS[16'h300F] = 8'h4D;
DFS[16'h3010] = 8'h61;
DFS[16'h3011] = 8'h74;
DFS[16'h3012] = 8'h68;
DFS[16'h3013] = 8'h65;
DFS[16'h3014] = 8'h72;
DFS[16'h3015] = 8'h20;
DFS[16'h3016] = 8'h28;
DFS[16'h3017] = 8'h31;
DFS[16'h3018] = 8'h39;
DFS[16'h3019] = 8'h20;
DFS[16'h301A] = 8'h4E;
DFS[16'h301B] = 8'h6F;
DFS[16'h301C] = 8'h76;
DFS[16'h301D] = 8'h20;
DFS[16'h301E] = 8'h32;
DFS[16'h301F] = 8'h30;
DFS[16'h3020] = 8'h30;
DFS[16'h3021] = 8'h38;
DFS[16'h3022] = 8'h29;
DFS[16'h3023] = 8'h00;
DFS[16'h3024] = 8'h4C;
DFS[16'h3025] = 8'hE7;
DFS[16'h3026] = 8'hFF;
DFS[16'h3027] = 8'hA2;
DFS[16'h3028] = 8'hFD;
DFS[16'h3029] = 8'h98;
DFS[16'h302A] = 8'h48;
DFS[16'h302B] = 8'hE8;
DFS[16'h302C] = 8'hE8;
DFS[16'h302D] = 8'h68;
DFS[16'h302E] = 8'h48;
DFS[16'h302F] = 8'hA8;
DFS[16'h3030] = 8'h20;
DFS[16'h3031] = 8'h6B;
DFS[16'h3032] = 8'hB0;
DFS[16'h3033] = 8'hE8;
DFS[16'h3034] = 8'hBD;
DFS[16'h3035] = 8'hF8;
DFS[16'h3036] = 8'hAE;
DFS[16'h3037] = 8'h30;
DFS[16'h3038] = 8'h28;
DFS[16'h3039] = 8'h86;
DFS[16'h303A] = 8'hB5;
DFS[16'h303B] = 8'hCA;
DFS[16'h303C] = 8'h88;
DFS[16'h303D] = 8'hE8;
DFS[16'h303E] = 8'hC8;
DFS[16'h303F] = 8'hBD;
DFS[16'h3040] = 8'hF8;
DFS[16'h3041] = 8'hAE;
DFS[16'h3042] = 8'h30;
DFS[16'h3043] = 8'h16;
DFS[16'h3044] = 8'h51;
DFS[16'h3045] = 8'hF2;
DFS[16'h3046] = 8'h29;
DFS[16'h3047] = 8'h5F;
DFS[16'h3048] = 8'hF0;
DFS[16'h3049] = 8'hF3;
DFS[16'h304A] = 8'hCA;
DFS[16'h304B] = 8'hE8;
DFS[16'h304C] = 8'hBD;
DFS[16'h304D] = 8'hF8;
DFS[16'h304E] = 8'hAE;
DFS[16'h304F] = 8'h10;
DFS[16'h3050] = 8'hFA;
DFS[16'h3051] = 8'hB1;
DFS[16'h3052] = 8'hF2;
DFS[16'h3053] = 8'hC9;
DFS[16'h3054] = 8'h2E;
DFS[16'h3055] = 8'hD0;
DFS[16'h3056] = 8'hD4;
DFS[16'h3057] = 8'hC8;
DFS[16'h3058] = 8'hB0;
DFS[16'h3059] = 8'h07;
DFS[16'h305A] = 8'hB1;
DFS[16'h305B] = 8'hF2;
DFS[16'h305C] = 8'h20;
DFS[16'h305D] = 8'hEE;
DFS[16'h305E] = 8'h82;
DFS[16'h305F] = 8'h90;
DFS[16'h3060] = 8'hCA;
DFS[16'h3061] = 8'h68;
DFS[16'h3062] = 8'hBD;
DFS[16'h3063] = 8'hF8;
DFS[16'h3064] = 8'hAE;
DFS[16'h3065] = 8'h48;
DFS[16'h3066] = 8'hBD;
DFS[16'h3067] = 8'hF9;
DFS[16'h3068] = 8'hAE;
DFS[16'h3069] = 8'h48;
DFS[16'h306A] = 8'h60;
DFS[16'h306B] = 8'hB1;
DFS[16'h306C] = 8'hF2;
DFS[16'h306D] = 8'hC9;
DFS[16'h306E] = 8'h0D;
DFS[16'h306F] = 8'hF0;
DFS[16'h3070] = 8'h08;
DFS[16'h3071] = 8'hC8;
DFS[16'h3072] = 8'hF0;
DFS[16'h3073] = 8'h07;
DFS[16'h3074] = 8'hC9;
DFS[16'h3075] = 8'h20;
DFS[16'h3076] = 8'hF0;
DFS[16'h3077] = 8'hF3;
DFS[16'h3078] = 8'h18;
DFS[16'h3079] = 8'h88;
DFS[16'h307A] = 8'h60;
DFS[16'h307B] = 8'h4C;
DFS[16'h307C] = 8'hB0;
DFS[16'h307D] = 8'hB2;
DFS[16'h307E] = 8'h98;
DFS[16'h307F] = 8'h48;
DFS[16'h3080] = 8'hA9;
DFS[16'h3081] = 8'h00;
DFS[16'h3082] = 8'h8D;
DFS[16'h3083] = 8'h55;
DFS[16'h3084] = 8'h0D;
DFS[16'h3085] = 8'h8D;
DFS[16'h3086] = 8'h56;
DFS[16'h3087] = 8'h0D;
DFS[16'h3088] = 8'h20;
DFS[16'h3089] = 8'h6B;
DFS[16'h308A] = 8'hB0;
DFS[16'h308B] = 8'hB0;
DFS[16'h308C] = 8'h62;
DFS[16'h308D] = 8'hB1;
DFS[16'h308E] = 8'hF2;
DFS[16'h308F] = 8'hC9;
DFS[16'h3090] = 8'h0D;
DFS[16'h3091] = 8'hF0;
DFS[16'h3092] = 8'h5C;
DFS[16'h3093] = 8'h38;
DFS[16'h3094] = 8'hE9;
DFS[16'h3095] = 8'h30;
DFS[16'h3096] = 8'h30;
DFS[16'h3097] = 8'h57;
DFS[16'h3098] = 8'hC9;
DFS[16'h3099] = 8'h0A;
DFS[16'h309A] = 8'hB0;
DFS[16'h309B] = 8'h53;
DFS[16'h309C] = 8'h48;
DFS[16'h309D] = 8'hAD;
DFS[16'h309E] = 8'h55;
DFS[16'h309F] = 8'h0D;
DFS[16'h30A0] = 8'h0A;
DFS[16'h30A1] = 8'h48;
DFS[16'h30A2] = 8'h2E;
DFS[16'h30A3] = 8'h56;
DFS[16'h30A4] = 8'h0D;
DFS[16'h30A5] = 8'hAE;
DFS[16'h30A6] = 8'h56;
DFS[16'h30A7] = 8'h0D;
DFS[16'h30A8] = 8'h0A;
DFS[16'h30A9] = 8'h2E;
DFS[16'h30AA] = 8'h56;
DFS[16'h30AB] = 8'h0D;
DFS[16'h30AC] = 8'h0A;
DFS[16'h30AD] = 8'h2E;
DFS[16'h30AE] = 8'h56;
DFS[16'h30AF] = 8'h0D;
DFS[16'h30B0] = 8'h8D;
DFS[16'h30B1] = 8'h55;
DFS[16'h30B2] = 8'h0D;
DFS[16'h30B3] = 8'h68;
DFS[16'h30B4] = 8'h6D;
DFS[16'h30B5] = 8'h55;
DFS[16'h30B6] = 8'h0D;
DFS[16'h30B7] = 8'h8D;
DFS[16'h30B8] = 8'h55;
DFS[16'h30B9] = 8'h0D;
DFS[16'h30BA] = 8'h8A;
DFS[16'h30BB] = 8'h6D;
DFS[16'h30BC] = 8'h56;
DFS[16'h30BD] = 8'h0D;
DFS[16'h30BE] = 8'hAA;
DFS[16'h30BF] = 8'h68;
DFS[16'h30C0] = 8'h6D;
DFS[16'h30C1] = 8'h55;
DFS[16'h30C2] = 8'h0D;
DFS[16'h30C3] = 8'h8D;
DFS[16'h30C4] = 8'h55;
DFS[16'h30C5] = 8'h0D;
DFS[16'h30C6] = 8'h8A;
DFS[16'h30C7] = 8'h69;
DFS[16'h30C8] = 8'h00;
DFS[16'h30C9] = 8'h8D;
DFS[16'h30CA] = 8'h56;
DFS[16'h30CB] = 8'h0D;
DFS[16'h30CC] = 8'hC9;
DFS[16'h30CD] = 8'h02;
DFS[16'h30CE] = 8'hB0;
DFS[16'h30CF] = 8'h1F;
DFS[16'h30D0] = 8'hC8;
DFS[16'h30D1] = 8'hF0;
DFS[16'h30D2] = 8'h1C;
DFS[16'h30D3] = 8'hB1;
DFS[16'h30D4] = 8'hF2;
DFS[16'h30D5] = 8'hC9;
DFS[16'h30D6] = 8'h0D;
DFS[16'h30D7] = 8'hF0;
DFS[16'h30D8] = 8'h04;
DFS[16'h30D9] = 8'hC9;
DFS[16'h30DA] = 8'h20;
DFS[16'h30DB] = 8'hD0;
DFS[16'h30DC] = 8'hB6;
DFS[16'h30DD] = 8'hAE;
DFS[16'h30DE] = 8'h55;
DFS[16'h30DF] = 8'h0D;
DFS[16'h30E0] = 8'hAD;
DFS[16'h30E1] = 8'h56;
DFS[16'h30E2] = 8'h0D;
DFS[16'h30E3] = 8'hF0;
DFS[16'h30E4] = 8'h04;
DFS[16'h30E5] = 8'hE8;
DFS[16'h30E6] = 8'hF0;
DFS[16'h30E7] = 8'h07;
DFS[16'h30E8] = 8'hCA;
DFS[16'h30E9] = 8'h68;
DFS[16'h30EA] = 8'hAD;
DFS[16'h30EB] = 8'h56;
DFS[16'h30EC] = 8'h0D;
DFS[16'h30ED] = 8'h18;
DFS[16'h30EE] = 8'h60;
DFS[16'h30EF] = 8'h68;
DFS[16'h30F0] = 8'hA8;
DFS[16'h30F1] = 8'hA9;
DFS[16'h30F2] = 8'h00;
DFS[16'h30F3] = 8'hAA;
DFS[16'h30F4] = 8'h38;
DFS[16'h30F5] = 8'h60;
DFS[16'h30F6] = 8'hA9;
DFS[16'h30F7] = 8'h0D;
DFS[16'h30F8] = 8'h8D;
DFS[16'h30F9] = 8'h5D;
DFS[16'h30FA] = 8'h0D;
DFS[16'h30FB] = 8'hA2;
DFS[16'h30FC] = 8'h00;
DFS[16'h30FD] = 8'h8E;
DFS[16'h30FE] = 8'h5E;
DFS[16'h30FF] = 8'h0D;
DFS[16'h3100] = 8'h20;
DFS[16'h3101] = 8'h6B;
DFS[16'h3102] = 8'hB0;
DFS[16'h3103] = 8'hB0;
DFS[16'h3104] = 8'h49;
DFS[16'h3105] = 8'hC9;
DFS[16'h3106] = 8'h22;
DFS[16'h3107] = 8'hD0;
DFS[16'h3108] = 8'h04;
DFS[16'h3109] = 8'hC8;
DFS[16'h310A] = 8'h8D;
DFS[16'h310B] = 8'h5D;
DFS[16'h310C] = 8'h0D;
DFS[16'h310D] = 8'hB1;
DFS[16'h310E] = 8'hF2;
DFS[16'h310F] = 8'hC9;
DFS[16'h3110] = 8'h0D;
DFS[16'h3111] = 8'hF0;
DFS[16'h3112] = 8'h2C;
DFS[16'h3113] = 8'hC9;
DFS[16'h3114] = 8'h20;
DFS[16'h3115] = 8'hD0;
DFS[16'h3116] = 8'h0B;
DFS[16'h3117] = 8'h90;
DFS[16'h3118] = 8'h52;
DFS[16'h3119] = 8'hAD;
DFS[16'h311A] = 8'h5D;
DFS[16'h311B] = 8'h0D;
DFS[16'h311C] = 8'hC9;
DFS[16'h311D] = 8'h22;
DFS[16'h311E] = 8'hD0;
DFS[16'h311F] = 8'h28;
DFS[16'h3120] = 8'hA9;
DFS[16'h3121] = 8'h20;
DFS[16'h3122] = 8'hC9;
DFS[16'h3123] = 8'h22;
DFS[16'h3124] = 8'hF0;
DFS[16'h3125] = 8'h19;
DFS[16'h3126] = 8'hC9;
DFS[16'h3127] = 8'h2A;
DFS[16'h3128] = 8'hF0;
DFS[16'h3129] = 8'h31;
DFS[16'h312A] = 8'hC9;
DFS[16'h312B] = 8'h61;
DFS[16'h312C] = 8'h90;
DFS[16'h312D] = 8'h06;
DFS[16'h312E] = 8'hC9;
DFS[16'h312F] = 8'h7B;
DFS[16'h3130] = 8'hB0;
DFS[16'h3131] = 8'h02;
DFS[16'h3132] = 8'h49;
DFS[16'h3133] = 8'h20;
DFS[16'h3134] = 8'h9D;
DFS[16'h3135] = 8'h5F;
DFS[16'h3136] = 8'h0D;
DFS[16'h3137] = 8'hC8;
DFS[16'h3138] = 8'hE8;
DFS[16'h3139] = 8'hE0;
DFS[16'h313A] = 8'h0C;
DFS[16'h313B] = 8'hD0;
DFS[16'h313C] = 8'hD0;
DFS[16'h313D] = 8'hB1;
DFS[16'h313E] = 8'hF2;
DFS[16'h313F] = 8'hCD;
DFS[16'h3140] = 8'h5D;
DFS[16'h3141] = 8'h0D;
DFS[16'h3142] = 8'hD0;
DFS[16'h3143] = 8'h27;
DFS[16'h3144] = 8'hC9;
DFS[16'h3145] = 8'h0D;
DFS[16'h3146] = 8'hF0;
DFS[16'h3147] = 8'h06;
DFS[16'h3148] = 8'hC8;
DFS[16'h3149] = 8'h20;
DFS[16'h314A] = 8'h6B;
DFS[16'h314B] = 8'hB0;
DFS[16'h314C] = 8'h90;
DFS[16'h314D] = 8'h1D;
DFS[16'h314E] = 8'h8E;
DFS[16'h314F] = 8'h5C;
DFS[16'h3150] = 8'h0D;
DFS[16'h3151] = 8'hE0;
DFS[16'h3152] = 8'h0C;
DFS[16'h3153] = 8'hF0;
DFS[16'h3154] = 8'h05;
DFS[16'h3155] = 8'hA9;
DFS[16'h3156] = 8'h00;
DFS[16'h3157] = 8'h9D;
DFS[16'h3158] = 8'h5F;
DFS[16'h3159] = 8'h0D;
DFS[16'h315A] = 8'h60;
DFS[16'h315B] = 8'h8D;
DFS[16'h315C] = 8'h5E;
DFS[16'h315D] = 8'h0D;
DFS[16'h315E] = 8'hAD;
DFS[16'h315F] = 8'h5D;
DFS[16'h3160] = 8'h0D;
DFS[16'h3161] = 8'hC9;
DFS[16'h3162] = 8'h0D;
DFS[16'h3163] = 8'hF0;
DFS[16'h3164] = 8'hE3;
DFS[16'h3165] = 8'hC8;
DFS[16'h3166] = 8'hB1;
DFS[16'h3167] = 8'hF2;
DFS[16'h3168] = 8'h4C;
DFS[16'h3169] = 8'h3F;
DFS[16'h316A] = 8'hB1;
DFS[16'h316B] = 8'h4C;
DFS[16'h316C] = 8'hB0;
DFS[16'h316D] = 8'hB2;
DFS[16'h316E] = 8'hA0;
DFS[16'h316F] = 8'h00;
DFS[16'h3170] = 8'hAE;
DFS[16'h3171] = 8'h5C;
DFS[16'h3172] = 8'h0D;
DFS[16'h3173] = 8'hF0;
DFS[16'h3174] = 8'h17;
DFS[16'h3175] = 8'hB1;
DFS[16'h3176] = 8'hF2;
DFS[16'h3177] = 8'hF0;
DFS[16'h3178] = 8'h25;
DFS[16'h3179] = 8'hC9;
DFS[16'h317A] = 8'h61;
DFS[16'h317B] = 8'h90;
DFS[16'h317C] = 8'h06;
DFS[16'h317D] = 8'hC9;
DFS[16'h317E] = 8'h7B;
DFS[16'h317F] = 8'hB0;
DFS[16'h3180] = 8'h02;
DFS[16'h3181] = 8'h49;
DFS[16'h3182] = 8'h20;
DFS[16'h3183] = 8'hD9;
DFS[16'h3184] = 8'h5F;
DFS[16'h3185] = 8'h0D;
DFS[16'h3186] = 8'hD0;
DFS[16'h3187] = 8'h16;
DFS[16'h3188] = 8'hC8;
DFS[16'h3189] = 8'hCA;
DFS[16'h318A] = 8'hD0;
DFS[16'h318B] = 8'hE9;
DFS[16'h318C] = 8'hB1;
DFS[16'h318D] = 8'hF2;
DFS[16'h318E] = 8'hF0;
DFS[16'h318F] = 8'h0C;
DFS[16'h3190] = 8'hAD;
DFS[16'h3191] = 8'h5C;
DFS[16'h3192] = 8'h0D;
DFS[16'h3193] = 8'hC9;
DFS[16'h3194] = 8'h0C;
DFS[16'h3195] = 8'hF0;
DFS[16'h3196] = 8'h05;
DFS[16'h3197] = 8'hAD;
DFS[16'h3198] = 8'h5E;
DFS[16'h3199] = 8'h0D;
DFS[16'h319A] = 8'hF0;
DFS[16'h319B] = 8'h02;
DFS[16'h319C] = 8'h18;
DFS[16'h319D] = 8'h60;
DFS[16'h319E] = 8'h38;
DFS[16'h319F] = 8'h60;
DFS[16'h31A0] = 8'hB0;
DFS[16'h31A1] = 8'h05;
DFS[16'h31A2] = 8'hA9;
DFS[16'h31A3] = 8'h20;
DFS[16'h31A4] = 8'h20;
DFS[16'h31A5] = 8'hEE;
DFS[16'h31A6] = 8'hFF;
DFS[16'h31A7] = 8'hA2;
DFS[16'h31A8] = 8'h20;
DFS[16'h31A9] = 8'hA0;
DFS[16'h31AA] = 8'h04;
DFS[16'h31AB] = 8'hAD;
DFS[16'h31AC] = 8'h56;
DFS[16'h31AD] = 8'h0D;
DFS[16'h31AE] = 8'h20;
DFS[16'h31AF] = 8'hE1;
DFS[16'h31B0] = 8'hB1;
DFS[16'h31B1] = 8'hAD;
DFS[16'h31B2] = 8'h55;
DFS[16'h31B3] = 8'h0D;
DFS[16'h31B4] = 8'h20;
DFS[16'h31B5] = 8'hE1;
DFS[16'h31B6] = 8'hB1;
DFS[16'h31B7] = 8'hA9;
DFS[16'h31B8] = 8'h20;
DFS[16'h31B9] = 8'h20;
DFS[16'h31BA] = 8'hEE;
DFS[16'h31BB] = 8'hFF;
DFS[16'h31BC] = 8'hA0;
DFS[16'h31BD] = 8'h00;
DFS[16'h31BE] = 8'hB1;
DFS[16'h31BF] = 8'hF2;
DFS[16'h31C0] = 8'hF0;
DFS[16'h31C1] = 8'h08;
DFS[16'h31C2] = 8'h20;
DFS[16'h31C3] = 8'hEE;
DFS[16'h31C4] = 8'hFF;
DFS[16'h31C5] = 8'hC8;
DFS[16'h31C6] = 8'hC0;
DFS[16'h31C7] = 8'h0C;
DFS[16'h31C8] = 8'hD0;
DFS[16'h31C9] = 8'hF4;
DFS[16'h31CA] = 8'hA9;
DFS[16'h31CB] = 8'h20;
DFS[16'h31CC] = 8'h20;
DFS[16'h31CD] = 8'hEE;
DFS[16'h31CE] = 8'hFF;
DFS[16'h31CF] = 8'hC8;
DFS[16'h31D0] = 8'hC0;
DFS[16'h31D1] = 8'h0D;
DFS[16'h31D2] = 8'hD0;
DFS[16'h31D3] = 8'hF8;
DFS[16'h31D4] = 8'hAA;
DFS[16'h31D5] = 8'hA0;
DFS[16'h31D6] = 8'h0F;
DFS[16'h31D7] = 8'hB1;
DFS[16'h31D8] = 8'hF2;
DFS[16'h31D9] = 8'hD0;
DFS[16'h31DA] = 8'h02;
DFS[16'h31DB] = 8'hA2;
DFS[16'h31DC] = 8'h50;
DFS[16'h31DD] = 8'h8A;
DFS[16'h31DE] = 8'h4C;
DFS[16'h31DF] = 8'hEE;
DFS[16'h31E0] = 8'hFF;
DFS[16'h31E1] = 8'h48;
DFS[16'h31E2] = 8'h4A;
DFS[16'h31E3] = 8'h4A;
DFS[16'h31E4] = 8'h4A;
DFS[16'h31E5] = 8'h4A;
DFS[16'h31E6] = 8'h20;
DFS[16'h31E7] = 8'hEA;
DFS[16'h31E8] = 8'hB1;
DFS[16'h31E9] = 8'h68;
DFS[16'h31EA] = 8'h29;
DFS[16'h31EB] = 8'h0F;
DFS[16'h31EC] = 8'hF0;
DFS[16'h31ED] = 8'h08;
DFS[16'h31EE] = 8'hA2;
DFS[16'h31EF] = 8'h30;
DFS[16'h31F0] = 8'h18;
DFS[16'h31F1] = 8'h69;
DFS[16'h31F2] = 8'h30;
DFS[16'h31F3] = 8'h4C;
DFS[16'h31F4] = 8'hEE;
DFS[16'h31F5] = 8'hFF;
DFS[16'h31F6] = 8'h88;
DFS[16'h31F7] = 8'hD0;
DFS[16'h31F8] = 8'h02;
DFS[16'h31F9] = 8'hA2;
DFS[16'h31FA] = 8'h30;
DFS[16'h31FB] = 8'h8A;
DFS[16'h31FC] = 8'h4C;
DFS[16'h31FD] = 8'hEE;
DFS[16'h31FE] = 8'hFF;
DFS[16'h31FF] = 8'hA2;
DFS[16'h3200] = 8'h00;
DFS[16'h3201] = 8'h68;
DFS[16'h3202] = 8'h85;
DFS[16'h3203] = 8'hA0;
DFS[16'h3204] = 8'h68;
DFS[16'h3205] = 8'h85;
DFS[16'h3206] = 8'hA1;
DFS[16'h3207] = 8'hA0;
DFS[16'h3208] = 8'h00;
DFS[16'h3209] = 8'hF0;
DFS[16'h320A] = 8'h07;
DFS[16'h320B] = 8'hB1;
DFS[16'h320C] = 8'hA0;
DFS[16'h320D] = 8'hF0;
DFS[16'h320E] = 8'h0B;
DFS[16'h320F] = 8'h20;
DFS[16'h3210] = 8'h21;
DFS[16'h3211] = 8'hB2;
DFS[16'h3212] = 8'hE6;
DFS[16'h3213] = 8'hA0;
DFS[16'h3214] = 8'hD0;
DFS[16'h3215] = 8'hF5;
DFS[16'h3216] = 8'hE6;
DFS[16'h3217] = 8'hA1;
DFS[16'h3218] = 8'hD0;
DFS[16'h3219] = 8'hF1;
DFS[16'h321A] = 8'hA5;
DFS[16'h321B] = 8'hA1;
DFS[16'h321C] = 8'h48;
DFS[16'h321D] = 8'hA5;
DFS[16'h321E] = 8'hA0;
DFS[16'h321F] = 8'h48;
DFS[16'h3220] = 8'h60;
DFS[16'h3221] = 8'hE0;
DFS[16'h3222] = 8'h00;
DFS[16'h3223] = 8'hD0;
DFS[16'h3224] = 8'h03;
DFS[16'h3225] = 8'h4C;
DFS[16'h3226] = 8'hEE;
DFS[16'h3227] = 8'hFF;
DFS[16'h3228] = 8'h9D;
DFS[16'h3229] = 8'h00;
DFS[16'h322A] = 8'h01;
DFS[16'h322B] = 8'hE8;
DFS[16'h322C] = 8'h60;
DFS[16'h322D] = 8'h08;
DFS[16'h322E] = 8'h10;
DFS[16'h322F] = 8'h1C;
DFS[16'h3230] = 8'h22;
DFS[16'h3231] = 8'h43;
DFS[16'h3232] = 8'h49;
DFS[16'h3233] = 8'h4F;
DFS[16'h3234] = 8'h58;
DFS[16'h3235] = 8'h28;
DFS[16'h3236] = 8'h3C;
DFS[16'h3237] = 8'h64;
DFS[16'h3238] = 8'h72;
DFS[16'h3239] = 8'h76;
DFS[16'h323A] = 8'h3E;
DFS[16'h323B] = 8'h29;
DFS[16'h323C] = 8'h00;
DFS[16'h323D] = 8'h3C;
DFS[16'h323E] = 8'h64;
DFS[16'h323F] = 8'h6E;
DFS[16'h3240] = 8'h6F;
DFS[16'h3241] = 8'h3E;
DFS[16'h3242] = 8'h2F;
DFS[16'h3243] = 8'h3C;
DFS[16'h3244] = 8'h64;
DFS[16'h3245] = 8'h73;
DFS[16'h3246] = 8'h70;
DFS[16'h3247] = 8'h3E;
DFS[16'h3248] = 8'h00;
DFS[16'h3249] = 8'h3C;
DFS[16'h324A] = 8'h64;
DFS[16'h324B] = 8'h6E;
DFS[16'h324C] = 8'h6F;
DFS[16'h324D] = 8'h3E;
DFS[16'h324E] = 8'h00;
DFS[16'h324F] = 8'h28;
DFS[16'h3250] = 8'h28;
DFS[16'h3251] = 8'h3C;
DFS[16'h3252] = 8'h66;
DFS[16'h3253] = 8'h72;
DFS[16'h3254] = 8'h6F;
DFS[16'h3255] = 8'h6D;
DFS[16'h3256] = 8'h20;
DFS[16'h3257] = 8'h64;
DFS[16'h3258] = 8'h6E;
DFS[16'h3259] = 8'h6F;
DFS[16'h325A] = 8'h3E;
DFS[16'h325B] = 8'h29;
DFS[16'h325C] = 8'h20;
DFS[16'h325D] = 8'h3C;
DFS[16'h325E] = 8'h74;
DFS[16'h325F] = 8'h6F;
DFS[16'h3260] = 8'h20;
DFS[16'h3261] = 8'h64;
DFS[16'h3262] = 8'h6E;
DFS[16'h3263] = 8'h6F;
DFS[16'h3264] = 8'h3E;
DFS[16'h3265] = 8'h29;
DFS[16'h3266] = 8'h20;
DFS[16'h3267] = 8'h28;
DFS[16'h3268] = 8'h3C;
DFS[16'h3269] = 8'h61;
DFS[16'h326A] = 8'h64;
DFS[16'h326B] = 8'h73;
DFS[16'h326C] = 8'h70;
DFS[16'h326D] = 8'h3E;
DFS[16'h326E] = 8'h29;
DFS[16'h326F] = 8'h00;
DFS[16'h3270] = 8'h3C;
DFS[16'h3271] = 8'h64;
DFS[16'h3272] = 8'h72;
DFS[16'h3273] = 8'h76;
DFS[16'h3274] = 8'h3E;
DFS[16'h3275] = 8'h00;
DFS[16'h3276] = 8'h3C;
DFS[16'h3277] = 8'h66;
DFS[16'h3278] = 8'h73;
DFS[16'h3279] = 8'h70;
DFS[16'h327A] = 8'h3E;
DFS[16'h327B] = 8'h00;
DFS[16'h327C] = 8'h28;
DFS[16'h327D] = 8'h3C;
DFS[16'h327E] = 8'h6D;
DFS[16'h327F] = 8'h6F;
DFS[16'h3280] = 8'h64;
DFS[16'h3281] = 8'h65;
DFS[16'h3282] = 8'h3E;
DFS[16'h3283] = 8'h29;
DFS[16'h3284] = 8'h00;
DFS[16'h3285] = 8'h28;
DFS[16'h3286] = 8'h3C;
DFS[16'h3287] = 8'h72;
DFS[16'h3288] = 8'h6F;
DFS[16'h3289] = 8'h6D;
DFS[16'h328A] = 8'h3E;
DFS[16'h328B] = 8'h29;
DFS[16'h328C] = 8'h00;
DFS[16'h328D] = 8'h48;
DFS[16'h328E] = 8'h4A;
DFS[16'h328F] = 8'h4A;
DFS[16'h3290] = 8'h4A;
DFS[16'h3291] = 8'h4A;
DFS[16'h3292] = 8'h20;
DFS[16'h3293] = 8'h98;
DFS[16'h3294] = 8'hB2;
DFS[16'h3295] = 8'h68;
DFS[16'h3296] = 8'h29;
DFS[16'h3297] = 8'h0F;
DFS[16'h3298] = 8'hA8;
DFS[16'h3299] = 8'hF0;
DFS[16'h329A] = 8'h14;
DFS[16'h329B] = 8'hA9;
DFS[16'h329C] = 8'h20;
DFS[16'h329D] = 8'h20;
DFS[16'h329E] = 8'h21;
DFS[16'h329F] = 8'hB2;
DFS[16'h32A0] = 8'hB9;
DFS[16'h32A1] = 8'h2C;
DFS[16'h32A2] = 8'hB2;
DFS[16'h32A3] = 8'hA8;
DFS[16'h32A4] = 8'hB9;
DFS[16'h32A5] = 8'h2D;
DFS[16'h32A6] = 8'hB2;
DFS[16'h32A7] = 8'hF0;
DFS[16'h32A8] = 8'h06;
DFS[16'h32A9] = 8'h20;
DFS[16'h32AA] = 8'h21;
DFS[16'h32AB] = 8'hB2;
DFS[16'h32AC] = 8'hC8;
DFS[16'h32AD] = 8'hD0;
DFS[16'h32AE] = 8'hF5;
DFS[16'h32AF] = 8'h60;
DFS[16'h32B0] = 8'hA2;
DFS[16'h32B1] = 8'h00;
DFS[16'h32B2] = 8'h8E;
DFS[16'h32B3] = 8'h00;
DFS[16'h32B4] = 8'h01;
DFS[16'h32B5] = 8'hE8;
DFS[16'h32B6] = 8'h20;
DFS[16'h32B7] = 8'h01;
DFS[16'h32B8] = 8'hB2;
DFS[16'h32B9] = 8'h1A;
DFS[16'h32BA] = 8'h53;
DFS[16'h32BB] = 8'h79;
DFS[16'h32BC] = 8'h6E;
DFS[16'h32BD] = 8'h74;
DFS[16'h32BE] = 8'h61;
DFS[16'h32BF] = 8'h78;
DFS[16'h32C0] = 8'h3A;
DFS[16'h32C1] = 8'h20;
DFS[16'h32C2] = 8'h00;
DFS[16'h32C3] = 8'hA4;
DFS[16'h32C4] = 8'hB5;
DFS[16'h32C5] = 8'hB9;
DFS[16'h32C6] = 8'hF8;
DFS[16'h32C7] = 8'hAE;
DFS[16'h32C8] = 8'h30;
DFS[16'h32C9] = 8'h06;
DFS[16'h32CA] = 8'h20;
DFS[16'h32CB] = 8'h21;
DFS[16'h32CC] = 8'hB2;
DFS[16'h32CD] = 8'hC8;
DFS[16'h32CE] = 8'hD0;
DFS[16'h32CF] = 8'hF5;
DFS[16'h32D0] = 8'hC8;
DFS[16'h32D1] = 8'hC8;
DFS[16'h32D2] = 8'hB9;
DFS[16'h32D3] = 8'hF8;
DFS[16'h32D4] = 8'hAE;
DFS[16'h32D5] = 8'hC8;
DFS[16'h32D6] = 8'h84;
DFS[16'h32D7] = 8'hB5;
DFS[16'h32D8] = 8'h20;
DFS[16'h32D9] = 8'h8D;
DFS[16'h32DA] = 8'hB2;
DFS[16'h32DB] = 8'hE0;
DFS[16'h32DC] = 8'h00;
DFS[16'h32DD] = 8'hF0;
DFS[16'h32DE] = 8'h08;
DFS[16'h32DF] = 8'hA9;
DFS[16'h32E0] = 8'h00;
DFS[16'h32E1] = 8'h9D;
DFS[16'h32E2] = 8'h00;
DFS[16'h32E3] = 8'h01;
DFS[16'h32E4] = 8'h4C;
DFS[16'h32E5] = 8'h00;
DFS[16'h32E6] = 8'h01;
DFS[16'h32E7] = 8'h60;
DFS[16'h32E8] = 8'h4C;
DFS[16'h32E9] = 8'hB0;
DFS[16'h32EA] = 8'hB2;
DFS[16'h32EB] = 8'h20;
DFS[16'h32EC] = 8'h6B;
DFS[16'h32ED] = 8'hB0;
DFS[16'h32EE] = 8'hB0;
DFS[16'h32EF] = 8'h17;
DFS[16'h32F0] = 8'h20;
DFS[16'h32F1] = 8'h7E;
DFS[16'h32F2] = 8'hB0;
DFS[16'h32F3] = 8'hB0;
DFS[16'h32F4] = 8'hBB;
DFS[16'h32F5] = 8'h48;
DFS[16'h32F6] = 8'h20;
DFS[16'h32F7] = 8'h6B;
DFS[16'h32F8] = 8'hB0;
DFS[16'h32F9] = 8'h68;
DFS[16'h32FA] = 8'h90;
DFS[16'h32FB] = 8'hB4;
DFS[16'h32FC] = 8'hD0;
DFS[16'h32FD] = 8'h26;
DFS[16'h32FE] = 8'h8A;
DFS[16'h32FF] = 8'h8D;
DFS[16'h3300] = 8'h5B;
DFS[16'h3301] = 8'h0D;
DFS[16'h3302] = 8'hC9;
DFS[16'h3303] = 8'h04;
DFS[16'h3304] = 8'hB0;
DFS[16'h3305] = 8'h1E;
DFS[16'h3306] = 8'h60;
DFS[16'h3307] = 8'hA5;
DFS[16'h3308] = 8'hCF;
DFS[16'h3309] = 8'h60;
DFS[16'h330A] = 8'h20;
DFS[16'h330B] = 8'h6B;
DFS[16'h330C] = 8'hB0;
DFS[16'h330D] = 8'hB0;
DFS[16'h330E] = 8'hA1;
DFS[16'h330F] = 8'h20;
DFS[16'h3310] = 8'h7E;
DFS[16'h3311] = 8'hB0;
DFS[16'h3312] = 8'hB0;
DFS[16'h3313] = 8'h9C;
DFS[16'h3314] = 8'h48;
DFS[16'h3315] = 8'h20;
DFS[16'h3316] = 8'h6B;
DFS[16'h3317] = 8'hB0;
DFS[16'h3318] = 8'h68;
DFS[16'h3319] = 8'h90;
DFS[16'h331A] = 8'h95;
DFS[16'h331B] = 8'h60;
DFS[16'h331C] = 8'h20;
DFS[16'h331D] = 8'h6B;
DFS[16'h331E] = 8'hB0;
DFS[16'h331F] = 8'hB0;
DFS[16'h3320] = 8'h8F;
DFS[16'h3321] = 8'h4C;
DFS[16'h3322] = 8'h75;
DFS[16'h3323] = 8'hB3;
DFS[16'h3324] = 8'h20;
DFS[16'h3325] = 8'h00;
DFS[16'h3326] = 8'hA0;
DFS[16'h3327] = 8'hCD;
DFS[16'h3328] = 8'h42;
DFS[16'h3329] = 8'h61;
DFS[16'h332A] = 8'h64;
DFS[16'h332B] = 8'h20;
DFS[16'h332C] = 8'h64;
DFS[16'h332D] = 8'h72;
DFS[16'h332E] = 8'h69;
DFS[16'h332F] = 8'h76;
DFS[16'h3330] = 8'h65;
DFS[16'h3331] = 8'h00;
DFS[16'h3332] = 8'h20;
DFS[16'h3333] = 8'h00;
DFS[16'h3334] = 8'hA0;
DFS[16'h3335] = 8'hD6;
DFS[16'h3336] = 8'h44;
DFS[16'h3337] = 8'h69;
DFS[16'h3338] = 8'h73;
DFS[16'h3339] = 8'h6B;
DFS[16'h333A] = 8'h20;
DFS[16'h333B] = 8'h6E;
DFS[16'h333C] = 8'h6F;
DFS[16'h333D] = 8'h74;
DFS[16'h333E] = 8'h20;
DFS[16'h333F] = 8'h66;
DFS[16'h3340] = 8'h6F;
DFS[16'h3341] = 8'h75;
DFS[16'h3342] = 8'h6E;
DFS[16'h3343] = 8'h64;
DFS[16'h3344] = 8'h00;
DFS[16'h3345] = 8'h20;
DFS[16'h3346] = 8'h6B;
DFS[16'h3347] = 8'hB0;
DFS[16'h3348] = 8'hB0;
DFS[16'h3349] = 8'h9E;
DFS[16'h334A] = 8'hA9;
DFS[16'h334B] = 8'hFF;
DFS[16'h334C] = 8'h20;
DFS[16'h334D] = 8'h5D;
DFS[16'h334E] = 8'hB3;
DFS[16'h334F] = 8'h08;
DFS[16'h3350] = 8'hE0;
DFS[16'h3351] = 8'h04;
DFS[16'h3352] = 8'hB0;
DFS[16'h3353] = 8'h33;
DFS[16'h3354] = 8'h28;
DFS[16'h3355] = 8'h60;
DFS[16'h3356] = 8'h20;
DFS[16'h3357] = 8'h6B;
DFS[16'h3358] = 8'hB0;
DFS[16'h3359] = 8'hB0;
DFS[16'h335A] = 8'h8D;
DFS[16'h335B] = 8'hA5;
DFS[16'h335C] = 8'hCF;
DFS[16'h335D] = 8'h8D;
DFS[16'h335E] = 8'h5B;
DFS[16'h335F] = 8'h0D;
DFS[16'h3360] = 8'h20;
DFS[16'h3361] = 8'h7E;
DFS[16'h3362] = 8'hB0;
DFS[16'h3363] = 8'hB0;
DFS[16'h3364] = 8'h26;
DFS[16'h3365] = 8'h48;
DFS[16'h3366] = 8'h20;
DFS[16'h3367] = 8'h6B;
DFS[16'h3368] = 8'hB0;
DFS[16'h3369] = 8'hB0;
DFS[16'h336A] = 8'h15;
DFS[16'h336B] = 8'h68;
DFS[16'h336C] = 8'hD0;
DFS[16'h336D] = 8'hB6;
DFS[16'h336E] = 8'hE0;
DFS[16'h336F] = 8'h04;
DFS[16'h3370] = 8'hB0;
DFS[16'h3371] = 8'hB2;
DFS[16'h3372] = 8'h8E;
DFS[16'h3373] = 8'h5B;
DFS[16'h3374] = 8'h0D;
DFS[16'h3375] = 8'h20;
DFS[16'h3376] = 8'h7E;
DFS[16'h3377] = 8'hB0;
DFS[16'h3378] = 8'hB0;
DFS[16'h3379] = 8'h11;
DFS[16'h337A] = 8'h48;
DFS[16'h337B] = 8'h20;
DFS[16'h337C] = 8'h6B;
DFS[16'h337D] = 8'hB0;
DFS[16'h337E] = 8'h90;
DFS[16'h337F] = 8'h07;
DFS[16'h3380] = 8'h68;
DFS[16'h3381] = 8'h6A;
DFS[16'h3382] = 8'h8A;
DFS[16'h3383] = 8'hAE;
DFS[16'h3384] = 8'h5B;
DFS[16'h3385] = 8'h0D;
DFS[16'h3386] = 8'h60;
DFS[16'h3387] = 8'h68;
DFS[16'h3388] = 8'h4C;
DFS[16'h3389] = 8'hB0;
DFS[16'h338A] = 8'hB2;
DFS[16'h338B] = 8'h20;
DFS[16'h338C] = 8'hF6;
DFS[16'h338D] = 8'hB0;
DFS[16'h338E] = 8'h20;
DFS[16'h338F] = 8'hBB;
DFS[16'h3390] = 8'hAD;
DFS[16'h3391] = 8'hAD;
DFS[16'h3392] = 8'h5C;
DFS[16'h3393] = 8'h0D;
DFS[16'h3394] = 8'hF0;
DFS[16'h3395] = 8'hF2;
DFS[16'h3396] = 8'hAD;
DFS[16'h3397] = 8'h5E;
DFS[16'h3398] = 8'h0D;
DFS[16'h3399] = 8'hD0;
DFS[16'h339A] = 8'hED;
DFS[16'h339B] = 8'hAD;
DFS[16'h339C] = 8'h54;
DFS[16'h339D] = 8'h0D;
DFS[16'h339E] = 8'h30;
DFS[16'h339F] = 8'h92;
DFS[16'h33A0] = 8'h20;
DFS[16'h33A1] = 8'h6E;
DFS[16'h33A2] = 8'hB1;
DFS[16'h33A3] = 8'h90;
DFS[16'h33A4] = 8'h06;
DFS[16'h33A5] = 8'h20;
DFS[16'h33A6] = 8'hE0;
DFS[16'h33A7] = 8'hAD;
DFS[16'h33A8] = 8'h4C;
DFS[16'h33A9] = 8'h9B;
DFS[16'h33AA] = 8'hB3;
DFS[16'h33AB] = 8'hAD;
DFS[16'h33AC] = 8'h54;
DFS[16'h33AD] = 8'h0D;
DFS[16'h33AE] = 8'h6A;
DFS[16'h33AF] = 8'hAD;
DFS[16'h33B0] = 8'h53;
DFS[16'h33B1] = 8'h0D;
DFS[16'h33B2] = 8'hAE;
DFS[16'h33B3] = 8'h5B;
DFS[16'h33B4] = 8'h0D;
DFS[16'h33B5] = 8'h60;
DFS[16'h33B6] = 8'h20;
DFS[16'h33B7] = 8'h1C;
DFS[16'h33B8] = 8'hB3;
DFS[16'h33B9] = 8'hA6;
DFS[16'h33BA] = 8'hCF;
DFS[16'h33BB] = 8'h20;
DFS[16'h33BC] = 8'h1B;
DFS[16'h33BD] = 8'hAC;
DFS[16'h33BE] = 8'h4C;
DFS[16'h33BF] = 8'h07;
DFS[16'h33C0] = 8'h94;
DFS[16'h33C1] = 8'h20;
DFS[16'h33C2] = 8'h56;
DFS[16'h33C3] = 8'hB3;
DFS[16'h33C4] = 8'h4C;
DFS[16'h33C5] = 8'h1B;
DFS[16'h33C6] = 8'hAC;
DFS[16'h33C7] = 8'hA9;
DFS[16'h33C8] = 8'h00;
DFS[16'h33C9] = 8'h8D;
DFS[16'h33CA] = 8'h57;
DFS[16'h33CB] = 8'h0D;
DFS[16'h33CC] = 8'h8D;
DFS[16'h33CD] = 8'h58;
DFS[16'h33CE] = 8'h0D;
DFS[16'h33CF] = 8'h20;
DFS[16'h33D0] = 8'h7E;
DFS[16'h33D1] = 8'hB0;
DFS[16'h33D2] = 8'hB0;
DFS[16'h33D3] = 8'h2D;
DFS[16'h33D4] = 8'h8E;
DFS[16'h33D5] = 8'h59;
DFS[16'h33D6] = 8'h0D;
DFS[16'h33D7] = 8'h8E;
DFS[16'h33D8] = 8'h53;
DFS[16'h33D9] = 8'h0D;
DFS[16'h33DA] = 8'h8D;
DFS[16'h33DB] = 8'h5A;
DFS[16'h33DC] = 8'h0D;
DFS[16'h33DD] = 8'h8D;
DFS[16'h33DE] = 8'h54;
DFS[16'h33DF] = 8'h0D;
DFS[16'h33E0] = 8'h20;
DFS[16'h33E1] = 8'h7E;
DFS[16'h33E2] = 8'hB0;
DFS[16'h33E3] = 8'hB0;
DFS[16'h33E4] = 8'h25;
DFS[16'h33E5] = 8'h8E;
DFS[16'h33E6] = 8'h59;
DFS[16'h33E7] = 8'h0D;
DFS[16'h33E8] = 8'h8D;
DFS[16'h33E9] = 8'h5A;
DFS[16'h33EA] = 8'h0D;
DFS[16'h33EB] = 8'hEC;
DFS[16'h33EC] = 8'h53;
DFS[16'h33ED] = 8'h0D;
DFS[16'h33EE] = 8'hED;
DFS[16'h33EF] = 8'h54;
DFS[16'h33F0] = 8'h0D;
DFS[16'h33F1] = 8'h10;
DFS[16'h33F2] = 8'h1F;
DFS[16'h33F3] = 8'h20;
DFS[16'h33F4] = 8'h00;
DFS[16'h33F5] = 8'hA0;
DFS[16'h33F6] = 8'hFF;
DFS[16'h33F7] = 8'h42;
DFS[16'h33F8] = 8'h61;
DFS[16'h33F9] = 8'h64;
DFS[16'h33FA] = 8'h20;
DFS[16'h33FB] = 8'h72;
DFS[16'h33FC] = 8'h61;
DFS[16'h33FD] = 8'h6E;
DFS[16'h33FE] = 8'h67;
DFS[16'h33FF] = 8'h65;
DFS[16'h3400] = 8'h00;
DFS[16'h3401] = 8'hA2;
DFS[16'h3402] = 8'hFE;
DFS[16'h3403] = 8'h8E;
DFS[16'h3404] = 8'h59;
DFS[16'h3405] = 8'h0D;
DFS[16'h3406] = 8'hE8;
DFS[16'h3407] = 8'h8E;
DFS[16'h3408] = 8'h5A;
DFS[16'h3409] = 8'h0D;
DFS[16'h340A] = 8'hA9;
DFS[16'h340B] = 8'h00;
DFS[16'h340C] = 8'h8D;
DFS[16'h340D] = 8'h53;
DFS[16'h340E] = 8'h0D;
DFS[16'h340F] = 8'h8D;
DFS[16'h3410] = 8'h54;
DFS[16'h3411] = 8'h0D;
DFS[16'h3412] = 8'hEE;
DFS[16'h3413] = 8'h59;
DFS[16'h3414] = 8'h0D;
DFS[16'h3415] = 8'hD0;
DFS[16'h3416] = 8'h03;
DFS[16'h3417] = 8'hEE;
DFS[16'h3418] = 8'h5A;
DFS[16'h3419] = 8'h0D;
DFS[16'h341A] = 8'h20;
DFS[16'h341B] = 8'hF6;
DFS[16'h341C] = 8'hB0;
DFS[16'h341D] = 8'hAD;
DFS[16'h341E] = 8'h54;
DFS[16'h341F] = 8'h0D;
DFS[16'h3420] = 8'h6A;
DFS[16'h3421] = 8'hAD;
DFS[16'h3422] = 8'h53;
DFS[16'h3423] = 8'h0D;
DFS[16'h3424] = 8'h20;
DFS[16'h3425] = 8'h85;
DFS[16'h3426] = 8'hAD;
DFS[16'h3427] = 8'hA2;
DFS[16'h3428] = 8'h00;
DFS[16'h3429] = 8'hAD;
DFS[16'h342A] = 8'h5C;
DFS[16'h342B] = 8'h0D;
DFS[16'h342C] = 8'hD0;
DFS[16'h342D] = 8'h04;
DFS[16'h342E] = 8'hCA;
DFS[16'h342F] = 8'h8E;
DFS[16'h3430] = 8'h5E;
DFS[16'h3431] = 8'h0D;
DFS[16'h3432] = 8'hAD;
DFS[16'h3433] = 8'h54;
DFS[16'h3434] = 8'h0D;
DFS[16'h3435] = 8'h30;
DFS[16'h3436] = 8'h33;
DFS[16'h3437] = 8'hAD;
DFS[16'h3438] = 8'h53;
DFS[16'h3439] = 8'h0D;
DFS[16'h343A] = 8'hCD;
DFS[16'h343B] = 8'h59;
DFS[16'h343C] = 8'h0D;
DFS[16'h343D] = 8'hAD;
DFS[16'h343E] = 8'h54;
DFS[16'h343F] = 8'h0D;
DFS[16'h3440] = 8'hED;
DFS[16'h3441] = 8'h5A;
DFS[16'h3442] = 8'h0D;
DFS[16'h3443] = 8'hB0;
DFS[16'h3444] = 8'h25;
DFS[16'h3445] = 8'h20;
DFS[16'h3446] = 8'h6E;
DFS[16'h3447] = 8'hB1;
DFS[16'h3448] = 8'hB0;
DFS[16'h3449] = 8'h16;
DFS[16'h344A] = 8'h20;
DFS[16'h344B] = 8'hA0;
DFS[16'h344C] = 8'hB1;
DFS[16'h344D] = 8'hF8;
DFS[16'h344E] = 8'h18;
DFS[16'h344F] = 8'hAD;
DFS[16'h3450] = 8'h57;
DFS[16'h3451] = 8'h0D;
DFS[16'h3452] = 8'h69;
DFS[16'h3453] = 8'h01;
DFS[16'h3454] = 8'h8D;
DFS[16'h3455] = 8'h57;
DFS[16'h3456] = 8'h0D;
DFS[16'h3457] = 8'hAD;
DFS[16'h3458] = 8'h58;
DFS[16'h3459] = 8'h0D;
DFS[16'h345A] = 8'h69;
DFS[16'h345B] = 8'h00;
DFS[16'h345C] = 8'h8D;
DFS[16'h345D] = 8'h58;
DFS[16'h345E] = 8'h0D;
DFS[16'h345F] = 8'hD8;
DFS[16'h3460] = 8'h24;
DFS[16'h3461] = 8'hFF;
DFS[16'h3462] = 8'h30;
DFS[16'h3463] = 8'h47;
DFS[16'h3464] = 8'h20;
DFS[16'h3465] = 8'hE0;
DFS[16'h3466] = 8'hAD;
DFS[16'h3467] = 8'h4C;
DFS[16'h3468] = 8'h32;
DFS[16'h3469] = 8'hB4;
DFS[16'h346A] = 8'hA9;
DFS[16'h346B] = 8'h86;
DFS[16'h346C] = 8'h20;
DFS[16'h346D] = 8'hF4;
DFS[16'h346E] = 8'hFF;
DFS[16'h346F] = 8'hE0;
DFS[16'h3470] = 8'h00;
DFS[16'h3471] = 8'hF0;
DFS[16'h3472] = 8'h03;
DFS[16'h3473] = 8'h20;
DFS[16'h3474] = 8'hE7;
DFS[16'h3475] = 8'hFF;
DFS[16'h3476] = 8'hAD;
DFS[16'h3477] = 8'h58;
DFS[16'h3478] = 8'h0D;
DFS[16'h3479] = 8'hA2;
DFS[16'h347A] = 8'h00;
DFS[16'h347B] = 8'hA0;
DFS[16'h347C] = 8'h04;
DFS[16'h347D] = 8'h20;
DFS[16'h347E] = 8'hE1;
DFS[16'h347F] = 8'hB1;
DFS[16'h3480] = 8'hAD;
DFS[16'h3481] = 8'h57;
DFS[16'h3482] = 8'h0D;
DFS[16'h3483] = 8'h20;
DFS[16'h3484] = 8'hE1;
DFS[16'h3485] = 8'hB1;
DFS[16'h3486] = 8'h20;
DFS[16'h3487] = 8'hFF;
DFS[16'h3488] = 8'hB1;
DFS[16'h3489] = 8'h20;
DFS[16'h348A] = 8'h64;
DFS[16'h348B] = 8'h69;
DFS[16'h348C] = 8'h73;
DFS[16'h348D] = 8'h6B;
DFS[16'h348E] = 8'h00;
DFS[16'h348F] = 8'hAD;
DFS[16'h3490] = 8'h58;
DFS[16'h3491] = 8'h0D;
DFS[16'h3492] = 8'hD0;
DFS[16'h3493] = 8'h05;
DFS[16'h3494] = 8'hCE;
DFS[16'h3495] = 8'h57;
DFS[16'h3496] = 8'h0D;
DFS[16'h3497] = 8'hF0;
DFS[16'h3498] = 8'h05;
DFS[16'h3499] = 8'hA9;
DFS[16'h349A] = 8'h73;
DFS[16'h349B] = 8'h20;
DFS[16'h349C] = 8'hEE;
DFS[16'h349D] = 8'hFF;
DFS[16'h349E] = 8'h20;
DFS[16'h349F] = 8'hFF;
DFS[16'h34A0] = 8'hB1;
DFS[16'h34A1] = 8'h20;
DFS[16'h34A2] = 8'h66;
DFS[16'h34A3] = 8'h6F;
DFS[16'h34A4] = 8'h75;
DFS[16'h34A5] = 8'h6E;
DFS[16'h34A6] = 8'h64;
DFS[16'h34A7] = 8'h00;
DFS[16'h34A8] = 8'h4C;
DFS[16'h34A9] = 8'hE7;
DFS[16'h34AA] = 8'hFF;
DFS[16'h34AB] = 8'h4C;
DFS[16'h34AC] = 8'h82;
DFS[16'h34AD] = 8'hA0;
DFS[16'h34AE] = 8'h4C;
DFS[16'h34AF] = 8'hB0;
DFS[16'h34B0] = 8'hB2;
DFS[16'h34B1] = 8'h20;
DFS[16'h34B2] = 8'h6B;
DFS[16'h34B3] = 8'hB0;
DFS[16'h34B4] = 8'h90;
DFS[16'h34B5] = 8'hF8;
DFS[16'h34B6] = 8'hA2;
DFS[16'h34B7] = 8'h00;
DFS[16'h34B8] = 8'h8E;
DFS[16'h34B9] = 8'h57;
DFS[16'h34BA] = 8'h0D;
DFS[16'h34BB] = 8'h8E;
DFS[16'h34BC] = 8'h58;
DFS[16'h34BD] = 8'h0D;
DFS[16'h34BE] = 8'h8E;
DFS[16'h34BF] = 8'h59;
DFS[16'h34C0] = 8'h0D;
DFS[16'h34C1] = 8'h8E;
DFS[16'h34C2] = 8'h5A;
DFS[16'h34C3] = 8'h0D;
DFS[16'h34C4] = 8'hA9;
DFS[16'h34C5] = 8'h80;
DFS[16'h34C6] = 8'h20;
DFS[16'h34C7] = 8'h9C;
DFS[16'h34C8] = 8'hAC;
DFS[16'h34C9] = 8'hA9;
DFS[16'h34CA] = 8'h10;
DFS[16'h34CB] = 8'h85;
DFS[16'h34CC] = 8'hF2;
DFS[16'h34CD] = 8'hA9;
DFS[16'h34CE] = 8'h0E;
DFS[16'h34CF] = 8'h85;
DFS[16'h34D0] = 8'hF3;
DFS[16'h34D1] = 8'hA0;
DFS[16'h34D2] = 8'h0F;
DFS[16'h34D3] = 8'hB1;
DFS[16'h34D4] = 8'hF2;
DFS[16'h34D5] = 8'hC9;
DFS[16'h34D6] = 8'hFF;
DFS[16'h34D7] = 8'hF0;
DFS[16'h34D8] = 8'h42;
DFS[16'h34D9] = 8'hF8;
DFS[16'h34DA] = 8'hA8;
DFS[16'h34DB] = 8'h10;
DFS[16'h34DC] = 8'h0E;
DFS[16'h34DD] = 8'h18;
DFS[16'h34DE] = 8'hAD;
DFS[16'h34DF] = 8'h57;
DFS[16'h34E0] = 8'h0D;
DFS[16'h34E1] = 8'h69;
DFS[16'h34E2] = 8'h01;
DFS[16'h34E3] = 8'h8D;
DFS[16'h34E4] = 8'h57;
DFS[16'h34E5] = 8'h0D;
DFS[16'h34E6] = 8'h90;
DFS[16'h34E7] = 8'h03;
DFS[16'h34E8] = 8'hEE;
DFS[16'h34E9] = 8'h58;
DFS[16'h34EA] = 8'h0D;
DFS[16'h34EB] = 8'h18;
DFS[16'h34EC] = 8'hAD;
DFS[16'h34ED] = 8'h59;
DFS[16'h34EE] = 8'h0D;
DFS[16'h34EF] = 8'h69;
DFS[16'h34F0] = 8'h01;
DFS[16'h34F1] = 8'h8D;
DFS[16'h34F2] = 8'h59;
DFS[16'h34F3] = 8'h0D;
DFS[16'h34F4] = 8'h90;
DFS[16'h34F5] = 8'h03;
DFS[16'h34F6] = 8'hEE;
DFS[16'h34F7] = 8'h5A;
DFS[16'h34F8] = 8'h0D;
DFS[16'h34F9] = 8'hD8;
DFS[16'h34FA] = 8'h18;
DFS[16'h34FB] = 8'hA5;
DFS[16'h34FC] = 8'hF2;
DFS[16'h34FD] = 8'h69;
DFS[16'h34FE] = 8'h10;
DFS[16'h34FF] = 8'h85;
DFS[16'h3500] = 8'hF2;
DFS[16'h3501] = 8'hD0;
DFS[16'h3502] = 8'hCE;
DFS[16'h3503] = 8'hA5;
DFS[16'h3504] = 8'hF3;
DFS[16'h3505] = 8'h49;
DFS[16'h3506] = 8'h01;
DFS[16'h3507] = 8'h85;
DFS[16'h3508] = 8'hF3;
DFS[16'h3509] = 8'h6A;
DFS[16'h350A] = 8'hB0;
DFS[16'h350B] = 8'hC5;
DFS[16'h350C] = 8'hAD;
DFS[16'h350D] = 8'h82;
DFS[16'h350E] = 8'h10;
DFS[16'h350F] = 8'h69;
DFS[16'h3510] = 8'h02;
DFS[16'h3511] = 8'hC9;
DFS[16'h3512] = 8'hA0;
DFS[16'h3513] = 8'hF0;
DFS[16'h3514] = 8'h06;
DFS[16'h3515] = 8'h20;
DFS[16'h3516] = 8'h9C;
DFS[16'h3517] = 8'hAC;
DFS[16'h3518] = 8'h4C;
DFS[16'h3519] = 8'hD1;
DFS[16'h351A] = 8'hB4;
DFS[16'h351B] = 8'hA0;
DFS[16'h351C] = 8'h04;
DFS[16'h351D] = 8'hA2;
DFS[16'h351E] = 8'h00;
DFS[16'h351F] = 8'hAD;
DFS[16'h3520] = 8'h58;
DFS[16'h3521] = 8'h0D;
DFS[16'h3522] = 8'h20;
DFS[16'h3523] = 8'hE1;
DFS[16'h3524] = 8'hB1;
DFS[16'h3525] = 8'hAD;
DFS[16'h3526] = 8'h57;
DFS[16'h3527] = 8'h0D;
DFS[16'h3528] = 8'h20;
DFS[16'h3529] = 8'hE1;
DFS[16'h352A] = 8'hB1;
DFS[16'h352B] = 8'h20;
DFS[16'h352C] = 8'hFF;
DFS[16'h352D] = 8'hB1;
DFS[16'h352E] = 8'h20;
DFS[16'h352F] = 8'h6F;
DFS[16'h3530] = 8'h66;
DFS[16'h3531] = 8'h20;
DFS[16'h3532] = 8'h00;
DFS[16'h3533] = 8'hA2;
DFS[16'h3534] = 8'h00;
DFS[16'h3535] = 8'hA0;
DFS[16'h3536] = 8'h04;
DFS[16'h3537] = 8'hAD;
DFS[16'h3538] = 8'h5A;
DFS[16'h3539] = 8'h0D;
DFS[16'h353A] = 8'h20;
DFS[16'h353B] = 8'hE1;
DFS[16'h353C] = 8'hB1;
DFS[16'h353D] = 8'hAD;
DFS[16'h353E] = 8'h59;
DFS[16'h353F] = 8'h0D;
DFS[16'h3540] = 8'h20;
DFS[16'h3541] = 8'hE1;
DFS[16'h3542] = 8'hB1;
DFS[16'h3543] = 8'h20;
DFS[16'h3544] = 8'hFF;
DFS[16'h3545] = 8'hB1;
DFS[16'h3546] = 8'h20;
DFS[16'h3547] = 8'h64;
DFS[16'h3548] = 8'h69;
DFS[16'h3549] = 8'h73;
DFS[16'h354A] = 8'h6B;
DFS[16'h354B] = 8'h00;
DFS[16'h354C] = 8'hAD;
DFS[16'h354D] = 8'h5A;
DFS[16'h354E] = 8'h0D;
DFS[16'h354F] = 8'hD0;
DFS[16'h3550] = 8'h07;
DFS[16'h3551] = 8'hAD;
DFS[16'h3552] = 8'h59;
DFS[16'h3553] = 8'h0D;
DFS[16'h3554] = 8'hC9;
DFS[16'h3555] = 8'h01;
DFS[16'h3556] = 8'hF0;
DFS[16'h3557] = 8'h05;
DFS[16'h3558] = 8'hA9;
DFS[16'h3559] = 8'h73;
DFS[16'h355A] = 8'h20;
DFS[16'h355B] = 8'hEE;
DFS[16'h355C] = 8'hFF;
DFS[16'h355D] = 8'h20;
DFS[16'h355E] = 8'hFF;
DFS[16'h355F] = 8'hB1;
DFS[16'h3560] = 8'h20;
DFS[16'h3561] = 8'h66;
DFS[16'h3562] = 8'h72;
DFS[16'h3563] = 8'h65;
DFS[16'h3564] = 8'h65;
DFS[16'h3565] = 8'h20;
DFS[16'h3566] = 8'h28;
DFS[16'h3567] = 8'h75;
DFS[16'h3568] = 8'h6E;
DFS[16'h3569] = 8'h66;
DFS[16'h356A] = 8'h6F;
DFS[16'h356B] = 8'h72;
DFS[16'h356C] = 8'h6D;
DFS[16'h356D] = 8'h61;
DFS[16'h356E] = 8'h74;
DFS[16'h356F] = 8'h74;
DFS[16'h3570] = 8'h65;
DFS[16'h3571] = 8'h64;
DFS[16'h3572] = 8'h29;
DFS[16'h3573] = 8'h00;
DFS[16'h3574] = 8'h4C;
DFS[16'h3575] = 8'hE7;
DFS[16'h3576] = 8'hFF;
DFS[16'h3577] = 8'h20;
DFS[16'h3578] = 8'hEB;
DFS[16'h3579] = 8'hB2;
DFS[16'h357A] = 8'hA2;
DFS[16'h357B] = 8'h04;
DFS[16'h357C] = 8'h8E;
DFS[16'h357D] = 8'h5B;
DFS[16'h357E] = 8'h0D;
DFS[16'h357F] = 8'hA2;
DFS[16'h3580] = 8'h00;
DFS[16'h3581] = 8'hB0;
DFS[16'h3582] = 8'h06;
DFS[16'h3583] = 8'hAA;
DFS[16'h3584] = 8'hE8;
DFS[16'h3585] = 8'h8E;
DFS[16'h3586] = 8'h5B;
DFS[16'h3587] = 8'h0D;
DFS[16'h3588] = 8'hCA;
DFS[16'h3589] = 8'h8A;
DFS[16'h358A] = 8'h48;
DFS[16'h358B] = 8'hA2;
DFS[16'h358C] = 8'h20;
DFS[16'h358D] = 8'hA0;
DFS[16'h358E] = 8'h02;
DFS[16'h358F] = 8'h20;
DFS[16'h3590] = 8'hE1;
DFS[16'h3591] = 8'hB1;
DFS[16'h3592] = 8'hA9;
DFS[16'h3593] = 8'h3A;
DFS[16'h3594] = 8'h20;
DFS[16'h3595] = 8'hEE;
DFS[16'h3596] = 8'hFF;
DFS[16'h3597] = 8'h68;
DFS[16'h3598] = 8'hAA;
DFS[16'h3599] = 8'h48;
DFS[16'h359A] = 8'hBD;
DFS[16'h359B] = 8'h10;
DFS[16'h359C] = 8'h0D;
DFS[16'h359D] = 8'h30;
DFS[16'h359E] = 8'h0F;
DFS[16'h359F] = 8'h6A;
DFS[16'h35A0] = 8'hBD;
DFS[16'h35A1] = 8'h0C;
DFS[16'h35A2] = 8'h0D;
DFS[16'h35A3] = 8'h20;
DFS[16'h35A4] = 8'h85;
DFS[16'h35A5] = 8'hAD;
DFS[16'h35A6] = 8'hC9;
DFS[16'h35A7] = 8'hFF;
DFS[16'h35A8] = 8'hF0;
DFS[16'h35A9] = 8'h04;
DFS[16'h35AA] = 8'h38;
DFS[16'h35AB] = 8'h20;
DFS[16'h35AC] = 8'hA0;
DFS[16'h35AD] = 8'hB1;
DFS[16'h35AE] = 8'h20;
DFS[16'h35AF] = 8'hE7;
DFS[16'h35B0] = 8'hFF;
DFS[16'h35B1] = 8'h68;
DFS[16'h35B2] = 8'hAA;
DFS[16'h35B3] = 8'hE8;
DFS[16'h35B4] = 8'hEC;
DFS[16'h35B5] = 8'h5B;
DFS[16'h35B6] = 8'h0D;
DFS[16'h35B7] = 8'h90;
DFS[16'h35B8] = 8'hD0;
DFS[16'h35B9] = 8'h60;
DFS[16'h35BA] = 8'h4C;
DFS[16'h35BB] = 8'hB0;
DFS[16'h35BC] = 8'hB2;
DFS[16'h35BD] = 8'hA9;
DFS[16'h35BE] = 8'h00;
DFS[16'h35BF] = 8'hF0;
DFS[16'h35C0] = 8'h02;
DFS[16'h35C1] = 8'hA9;
DFS[16'h35C2] = 8'h0F;
DFS[16'h35C3] = 8'h48;
DFS[16'h35C4] = 8'h20;
DFS[16'h35C5] = 8'h1C;
DFS[16'h35C6] = 8'hB3;
DFS[16'h35C7] = 8'h20;
DFS[16'h35C8] = 8'hCD;
DFS[16'h35C9] = 8'hAB;
DFS[16'h35CA] = 8'h30;
DFS[16'h35CB] = 8'h0E;
DFS[16'h35CC] = 8'h68;
DFS[16'h35CD] = 8'hB0;
DFS[16'h35CE] = 8'h05;
DFS[16'h35CF] = 8'h99;
DFS[16'h35D0] = 8'h00;
DFS[16'h35D1] = 8'h0E;
DFS[16'h35D2] = 8'h90;
DFS[16'h35D3] = 8'h03;
DFS[16'h35D4] = 8'h99;
DFS[16'h35D5] = 8'h00;
DFS[16'h35D6] = 8'h0F;
DFS[16'h35D7] = 8'h4C;
DFS[16'h35D8] = 8'hCD;
DFS[16'h35D9] = 8'hAC;
DFS[16'h35DA] = 8'hC9;
DFS[16'h35DB] = 8'hFF;
DFS[16'h35DC] = 8'hF0;
DFS[16'h35DD] = 8'h03;
DFS[16'h35DE] = 8'h4C;
DFS[16'h35DF] = 8'h65;
DFS[16'h35E0] = 8'hAC;
DFS[16'h35E1] = 8'h4C;
DFS[16'h35E2] = 8'h4B;
DFS[16'h35E3] = 8'hAC;
DFS[16'h35E4] = 8'h20;
DFS[16'h35E5] = 8'hBD;
DFS[16'h35E6] = 8'h9B;
DFS[16'h35E7] = 8'h20;
DFS[16'h35E8] = 8'h0A;
DFS[16'h35E9] = 8'hB3;
DFS[16'h35EA] = 8'h6A;
DFS[16'h35EB] = 8'h08;
DFS[16'h35EC] = 8'h8A;
DFS[16'h35ED] = 8'h48;
DFS[16'h35EE] = 8'h20;
DFS[16'h35EF] = 8'hCD;
DFS[16'h35F0] = 8'hAB;
DFS[16'h35F1] = 8'h30;
DFS[16'h35F2] = 8'hE7;
DFS[16'h35F3] = 8'h68;
DFS[16'h35F4] = 8'h28;
DFS[16'h35F5] = 8'h20;
DFS[16'h35F6] = 8'h85;
DFS[16'h35F7] = 8'hAD;
DFS[16'h35F8] = 8'h20;
DFS[16'h35F9] = 8'hFF;
DFS[16'h35FA] = 8'hB1;
DFS[16'h35FB] = 8'h4B;
DFS[16'h35FC] = 8'h69;
DFS[16'h35FD] = 8'h6C;
DFS[16'h35FE] = 8'h6C;
DFS[16'h35FF] = 8'h00;
DFS[16'h3600] = 8'h38;
DFS[16'h3601] = 8'h20;
DFS[16'h3602] = 8'hA0;
DFS[16'h3603] = 8'hB1;
DFS[16'h3604] = 8'h20;
DFS[16'h3605] = 8'hFF;
DFS[16'h3606] = 8'hB1;
DFS[16'h3607] = 8'h20;
DFS[16'h3608] = 8'h3A;
DFS[16'h3609] = 8'h20;
DFS[16'h360A] = 8'h00;
DFS[16'h360B] = 8'h20;
DFS[16'h360C] = 8'h9E;
DFS[16'h360D] = 8'h9C;
DFS[16'h360E] = 8'h08;
DFS[16'h360F] = 8'h20;
DFS[16'h3610] = 8'hE7;
DFS[16'h3611] = 8'hFF;
DFS[16'h3612] = 8'h28;
DFS[16'h3613] = 8'hD0;
DFS[16'h3614] = 8'h09;
DFS[16'h3615] = 8'hA0;
DFS[16'h3616] = 8'h0F;
DFS[16'h3617] = 8'hA9;
DFS[16'h3618] = 8'hF0;
DFS[16'h3619] = 8'h91;
DFS[16'h361A] = 8'hF2;
DFS[16'h361B] = 8'h4C;
DFS[16'h361C] = 8'hCD;
DFS[16'h361D] = 8'hAC;
DFS[16'h361E] = 8'h60;
DFS[16'h361F] = 8'hA9;
DFS[16'h3620] = 8'h00;
DFS[16'h3621] = 8'h20;
DFS[16'h3622] = 8'h29;
DFS[16'h3623] = 8'hB6;
DFS[16'h3624] = 8'h4C;
DFS[16'h3625] = 8'h6F;
DFS[16'h3626] = 8'hAB;
DFS[16'h3627] = 8'hA9;
DFS[16'h3628] = 8'h01;
DFS[16'h3629] = 8'h8D;
DFS[16'h362A] = 8'h5F;
DFS[16'h362B] = 8'h0D;
DFS[16'h362C] = 8'h20;
DFS[16'h362D] = 8'h0A;
DFS[16'h362E] = 8'hB3;
DFS[16'h362F] = 8'h6A;
DFS[16'h3630] = 8'h08;
DFS[16'h3631] = 8'h8A;
DFS[16'h3632] = 8'h48;
DFS[16'h3633] = 8'h20;
DFS[16'h3634] = 8'hCD;
DFS[16'h3635] = 8'hAB;
DFS[16'h3636] = 8'h10;
DFS[16'h3637] = 8'h26;
DFS[16'h3638] = 8'hAA;
DFS[16'h3639] = 8'hE8;
DFS[16'h363A] = 8'hF0;
DFS[16'h363B] = 8'h3D;
DFS[16'h363C] = 8'h98;
DFS[16'h363D] = 8'h29;
DFS[16'h363E] = 8'hF0;
DFS[16'h363F] = 8'h85;
DFS[16'h3640] = 8'hF2;
DFS[16'h3641] = 8'hA0;
DFS[16'h3642] = 8'h0E;
DFS[16'h3643] = 8'h90;
DFS[16'h3644] = 8'h01;
DFS[16'h3645] = 8'hC8;
DFS[16'h3646] = 8'h84;
DFS[16'h3647] = 8'hF3;
DFS[16'h3648] = 8'hA0;
DFS[16'h3649] = 8'h0F;
DFS[16'h364A] = 8'h98;
DFS[16'h364B] = 8'h91;
DFS[16'h364C] = 8'hF2;
DFS[16'h364D] = 8'hAD;
DFS[16'h364E] = 8'h5F;
DFS[16'h364F] = 8'h0D;
DFS[16'h3650] = 8'hD0;
DFS[16'h3651] = 8'h06;
DFS[16'h3652] = 8'h88;
DFS[16'h3653] = 8'h91;
DFS[16'h3654] = 8'hF2;
DFS[16'h3655] = 8'h88;
DFS[16'h3656] = 8'h10;
DFS[16'h3657] = 8'hFB;
DFS[16'h3658] = 8'h20;
DFS[16'h3659] = 8'hCD;
DFS[16'h365A] = 8'hAC;
DFS[16'h365B] = 8'h68;
DFS[16'h365C] = 8'h28;
DFS[16'h365D] = 8'h60;
DFS[16'h365E] = 8'h20;
DFS[16'h365F] = 8'h00;
DFS[16'h3660] = 8'hA0;
DFS[16'h3661] = 8'hFF;
DFS[16'h3662] = 8'h44;
DFS[16'h3663] = 8'h69;
DFS[16'h3664] = 8'h73;
DFS[16'h3665] = 8'h6B;
DFS[16'h3666] = 8'h20;
DFS[16'h3667] = 8'h61;
DFS[16'h3668] = 8'h6C;
DFS[16'h3669] = 8'h72;
DFS[16'h366A] = 8'h65;
DFS[16'h366B] = 8'h61;
DFS[16'h366C] = 8'h64;
DFS[16'h366D] = 8'h79;
DFS[16'h366E] = 8'h20;
DFS[16'h366F] = 8'h66;
DFS[16'h3670] = 8'h6F;
DFS[16'h3671] = 8'h72;
DFS[16'h3672] = 8'h6D;
DFS[16'h3673] = 8'h61;
DFS[16'h3674] = 8'h74;
DFS[16'h3675] = 8'h74;
DFS[16'h3676] = 8'h65;
DFS[16'h3677] = 8'h64;
DFS[16'h3678] = 8'h00;
DFS[16'h3679] = 8'h4C;
DFS[16'h367A] = 8'h4B;
DFS[16'h367B] = 8'hAC;
DFS[16'h367C] = 8'h20;
DFS[16'h367D] = 8'hEB;
DFS[16'h367E] = 8'hB2;
DFS[16'h367F] = 8'h8D;
DFS[16'h3680] = 8'h5B;
DFS[16'h3681] = 8'h0D;
DFS[16'h3682] = 8'h20;
DFS[16'h3683] = 8'hE0;
DFS[16'h3684] = 8'hB6;
DFS[16'h3685] = 8'h08;
DFS[16'h3686] = 8'h48;
DFS[16'h3687] = 8'hA9;
DFS[16'h3688] = 8'h0F;
DFS[16'h3689] = 8'h91;
DFS[16'h368A] = 8'hF2;
DFS[16'h368B] = 8'h88;
DFS[16'h368C] = 8'hA9;
DFS[16'h368D] = 8'h00;
DFS[16'h368E] = 8'h91;
DFS[16'h368F] = 8'hF2;
DFS[16'h3690] = 8'h88;
DFS[16'h3691] = 8'h10;
DFS[16'h3692] = 8'hFB;
DFS[16'h3693] = 8'h20;
DFS[16'h3694] = 8'hB8;
DFS[16'h3695] = 8'hAC;
DFS[16'h3696] = 8'h68;
DFS[16'h3697] = 8'h28;
DFS[16'h3698] = 8'h08;
DFS[16'h3699] = 8'h48;
DFS[16'h369A] = 8'h20;
DFS[16'h369B] = 8'h6F;
DFS[16'h369C] = 8'hAB;
DFS[16'h369D] = 8'h68;
DFS[16'h369E] = 8'h28;
DFS[16'h369F] = 8'h08;
DFS[16'h36A0] = 8'h48;
DFS[16'h36A1] = 8'hAE;
DFS[16'h36A2] = 8'h5B;
DFS[16'h36A3] = 8'h0D;
DFS[16'h36A4] = 8'h20;
DFS[16'h36A5] = 8'h1B;
DFS[16'h36A6] = 8'hAC;
DFS[16'h36A7] = 8'h20;
DFS[16'h36A8] = 8'hFF;
DFS[16'h36A9] = 8'hB1;
DFS[16'h36AA] = 8'h44;
DFS[16'h36AB] = 8'h69;
DFS[16'h36AC] = 8'h73;
DFS[16'h36AD] = 8'h6B;
DFS[16'h36AE] = 8'h20;
DFS[16'h36AF] = 8'h00;
DFS[16'h36B0] = 8'h68;
DFS[16'h36B1] = 8'h28;
DFS[16'h36B2] = 8'h20;
DFS[16'h36B3] = 8'hCD;
DFS[16'h36B4] = 8'hA9;
DFS[16'h36B5] = 8'h8E;
DFS[16'h36B6] = 8'h55;
DFS[16'h36B7] = 8'h0D;
DFS[16'h36B8] = 8'hA2;
DFS[16'h36B9] = 8'h00;
DFS[16'h36BA] = 8'hA0;
DFS[16'h36BB] = 8'h04;
DFS[16'h36BC] = 8'h20;
DFS[16'h36BD] = 8'hE1;
DFS[16'h36BE] = 8'hB1;
DFS[16'h36BF] = 8'hAD;
DFS[16'h36C0] = 8'h55;
DFS[16'h36C1] = 8'h0D;
DFS[16'h36C2] = 8'h20;
DFS[16'h36C3] = 8'hE1;
DFS[16'h36C4] = 8'hB1;
DFS[16'h36C5] = 8'h20;
DFS[16'h36C6] = 8'hFF;
DFS[16'h36C7] = 8'hB1;
DFS[16'h36C8] = 8'h20;
DFS[16'h36C9] = 8'h69;
DFS[16'h36CA] = 8'h6E;
DFS[16'h36CB] = 8'h20;
DFS[16'h36CC] = 8'h64;
DFS[16'h36CD] = 8'h72;
DFS[16'h36CE] = 8'h69;
DFS[16'h36CF] = 8'h76;
DFS[16'h36D0] = 8'h65;
DFS[16'h36D1] = 8'h20;
DFS[16'h36D2] = 8'h00;
DFS[16'h36D3] = 8'hAD;
DFS[16'h36D4] = 8'h5B;
DFS[16'h36D5] = 8'h0D;
DFS[16'h36D6] = 8'hA2;
DFS[16'h36D7] = 8'h00;
DFS[16'h36D8] = 8'hA0;
DFS[16'h36D9] = 8'h02;
DFS[16'h36DA] = 8'h20;
DFS[16'h36DB] = 8'hE1;
DFS[16'h36DC] = 8'hB1;
DFS[16'h36DD] = 8'h4C;
DFS[16'h36DE] = 8'hE7;
DFS[16'h36DF] = 8'hFF;
DFS[16'h36E0] = 8'hA9;
DFS[16'h36E1] = 8'h10;
DFS[16'h36E2] = 8'h85;
DFS[16'h36E3] = 8'hF2;
DFS[16'h36E4] = 8'hA9;
DFS[16'h36E5] = 8'h0E;
DFS[16'h36E6] = 8'h85;
DFS[16'h36E7] = 8'hF3;
DFS[16'h36E8] = 8'hA9;
DFS[16'h36E9] = 8'h80;
DFS[16'h36EA] = 8'h8D;
DFS[16'h36EB] = 8'h52;
DFS[16'h36EC] = 8'h0D;
DFS[16'h36ED] = 8'h20;
DFS[16'h36EE] = 8'hA1;
DFS[16'h36EF] = 8'hAC;
DFS[16'h36F0] = 8'hA9;
DFS[16'h36F1] = 8'h00;
DFS[16'h36F2] = 8'h8D;
DFS[16'h36F3] = 8'h53;
DFS[16'h36F4] = 8'h0D;
DFS[16'h36F5] = 8'h8D;
DFS[16'h36F6] = 8'h54;
DFS[16'h36F7] = 8'h0D;
DFS[16'h36F8] = 8'hA0;
DFS[16'h36F9] = 8'h0F;
DFS[16'h36FA] = 8'hB1;
DFS[16'h36FB] = 8'hF2;
DFS[16'h36FC] = 8'h10;
DFS[16'h36FD] = 8'h0C;
DFS[16'h36FE] = 8'hC9;
DFS[16'h36FF] = 8'hFF;
DFS[16'h3700] = 8'hF0;
DFS[16'h3701] = 8'h36;
DFS[16'h3702] = 8'hAD;
DFS[16'h3703] = 8'h54;
DFS[16'h3704] = 8'h0D;
DFS[16'h3705] = 8'h6A;
DFS[16'h3706] = 8'hAD;
DFS[16'h3707] = 8'h53;
DFS[16'h3708] = 8'h0D;
DFS[16'h3709] = 8'h60;
DFS[16'h370A] = 8'hEE;
DFS[16'h370B] = 8'h53;
DFS[16'h370C] = 8'h0D;
DFS[16'h370D] = 8'hD0;
DFS[16'h370E] = 8'h03;
DFS[16'h370F] = 8'hEE;
DFS[16'h3710] = 8'h54;
DFS[16'h3711] = 8'h0D;
DFS[16'h3712] = 8'h18;
DFS[16'h3713] = 8'hA5;
DFS[16'h3714] = 8'hF2;
DFS[16'h3715] = 8'h69;
DFS[16'h3716] = 8'h10;
DFS[16'h3717] = 8'h85;
DFS[16'h3718] = 8'hF2;
DFS[16'h3719] = 8'hD0;
DFS[16'h371A] = 8'hDF;
DFS[16'h371B] = 8'hA5;
DFS[16'h371C] = 8'hF3;
DFS[16'h371D] = 8'h49;
DFS[16'h371E] = 8'h01;
DFS[16'h371F] = 8'h85;
DFS[16'h3720] = 8'hF3;
DFS[16'h3721] = 8'h29;
DFS[16'h3722] = 8'h01;
DFS[16'h3723] = 8'hD0;
DFS[16'h3724] = 8'hD5;
DFS[16'h3725] = 8'h18;
DFS[16'h3726] = 8'hAD;
DFS[16'h3727] = 8'h52;
DFS[16'h3728] = 8'h0D;
DFS[16'h3729] = 8'h69;
DFS[16'h372A] = 8'h02;
DFS[16'h372B] = 8'hC9;
DFS[16'h372C] = 8'hA0;
DFS[16'h372D] = 8'hF0;
DFS[16'h372E] = 8'h09;
DFS[16'h372F] = 8'h8D;
DFS[16'h3730] = 8'h52;
DFS[16'h3731] = 8'h0D;
DFS[16'h3732] = 8'h20;
DFS[16'h3733] = 8'hA1;
DFS[16'h3734] = 8'hAC;
DFS[16'h3735] = 8'h4C;
DFS[16'h3736] = 8'hF8;
DFS[16'h3737] = 8'hB6;
DFS[16'h3738] = 8'h20;
DFS[16'h3739] = 8'h00;
DFS[16'h373A] = 8'hA0;
DFS[16'h373B] = 8'hFF;
DFS[16'h373C] = 8'h4E;
DFS[16'h373D] = 8'h6F;
DFS[16'h373E] = 8'h20;
DFS[16'h373F] = 8'h66;
DFS[16'h3740] = 8'h72;
DFS[16'h3741] = 8'h65;
DFS[16'h3742] = 8'h65;
DFS[16'h3743] = 8'h20;
DFS[16'h3744] = 8'h64;
DFS[16'h3745] = 8'h69;
DFS[16'h3746] = 8'h73;
DFS[16'h3747] = 8'h6B;
DFS[16'h3748] = 8'h73;
DFS[16'h3749] = 8'h00;
DFS[16'h374A] = 8'h20;
DFS[16'h374B] = 8'h45;
DFS[16'h374C] = 8'hB3;
DFS[16'h374D] = 8'h08;
DFS[16'h374E] = 8'h48;
DFS[16'h374F] = 8'h8A;
DFS[16'h3750] = 8'h48;
DFS[16'h3751] = 8'hA9;
DFS[16'h3752] = 8'h80;
DFS[16'h3753] = 8'h20;
DFS[16'h3754] = 8'hA1;
DFS[16'h3755] = 8'hAC;
DFS[16'h3756] = 8'h68;
DFS[16'h3757] = 8'hAA;
DFS[16'h3758] = 8'h68;
DFS[16'h3759] = 8'h9D;
DFS[16'h375A] = 8'h00;
DFS[16'h375B] = 8'h0E;
DFS[16'h375C] = 8'h68;
DFS[16'h375D] = 8'h29;
DFS[16'h375E] = 8'h01;
DFS[16'h375F] = 8'h9D;
DFS[16'h3760] = 8'h04;
DFS[16'h3761] = 8'h0E;
DFS[16'h3762] = 8'h4C;
DFS[16'h3763] = 8'hB8;
DFS[16'h3764] = 8'hAC;
DFS[16'h3765] = 8'h20;
DFS[16'h3766] = 8'h6B;
DFS[16'h3767] = 8'hB0;
DFS[16'h3768] = 8'hA2;
DFS[16'h3769] = 8'h00;
DFS[16'h376A] = 8'hB0;
DFS[16'h376B] = 8'h0B;
DFS[16'h376C] = 8'h20;
DFS[16'h376D] = 8'h7E;
DFS[16'h376E] = 8'hB0;
DFS[16'h376F] = 8'hB0;
DFS[16'h3770] = 8'h16;
DFS[16'h3771] = 8'hC9;
DFS[16'h3772] = 8'h00;
DFS[16'h3773] = 8'hF0;
DFS[16'h3774] = 8'h02;
DFS[16'h3775] = 8'hA2;
DFS[16'h3776] = 8'h01;
DFS[16'h3777] = 8'h8E;
DFS[16'h3778] = 8'h04;
DFS[16'h3779] = 8'h0D;
DFS[16'h377A] = 8'h20;
DFS[16'h377B] = 8'hE2;
DFS[16'h377C] = 8'h8D;
DFS[16'h377D] = 8'hA2;
DFS[16'h377E] = 8'hFF;
DFS[16'h377F] = 8'hA9;
DFS[16'h3780] = 8'h61;
DFS[16'h3781] = 8'h8D;
DFS[16'h3782] = 8'h52;
DFS[16'h3783] = 8'h0D;
DFS[16'h3784] = 8'h4C;
DFS[16'h3785] = 8'h17;
DFS[16'h3786] = 8'hAD;
DFS[16'h3787] = 8'h20;
DFS[16'h3788] = 8'h00;
DFS[16'h3789] = 8'hA0;
DFS[16'h378A] = 8'hFF;
DFS[16'h378B] = 8'h42;
DFS[16'h378C] = 8'h61;
DFS[16'h378D] = 8'h64;
DFS[16'h378E] = 8'h20;
DFS[16'h378F] = 8'h64;
DFS[16'h3790] = 8'h72;
DFS[16'h3791] = 8'h69;
DFS[16'h3792] = 8'h76;
DFS[16'h3793] = 8'h65;
DFS[16'h3794] = 8'h72;
DFS[16'h3795] = 8'h20;
DFS[16'h3796] = 8'h6D;
DFS[16'h3797] = 8'h6F;
DFS[16'h3798] = 8'h64;
DFS[16'h3799] = 8'h65;
DFS[16'h379A] = 8'h00;
DFS[16'h379B] = 8'hA2;
DFS[16'h379C] = 8'h1E;
DFS[16'h379D] = 8'hBC;
DFS[16'h379E] = 8'h02;
DFS[16'h379F] = 8'h0D;
DFS[16'h37A0] = 8'hBD;
DFS[16'h37A1] = 8'h21;
DFS[16'h37A2] = 8'h0D;
DFS[16'h37A3] = 8'h9D;
DFS[16'h37A4] = 8'h02;
DFS[16'h37A5] = 8'h0D;
DFS[16'h37A6] = 8'h98;
DFS[16'h37A7] = 8'h9D;
DFS[16'h37A8] = 8'h21;
DFS[16'h37A9] = 8'h0D;
DFS[16'h37AA] = 8'hCA;
DFS[16'h37AB] = 8'h10;
DFS[16'h37AC] = 8'hF0;
DFS[16'h37AD] = 8'h8E;
DFS[16'h37AE] = 8'h82;
DFS[16'h37AF] = 8'h10;
DFS[16'h37B0] = 8'h60;
DFS[16'h37B1] = 8'hA9;
DFS[16'h37B2] = 8'h00;
DFS[16'h37B3] = 8'h85;
DFS[16'h37B4] = 8'hA6;
DFS[16'h37B5] = 8'h20;
DFS[16'h37B6] = 8'hC2;
DFS[16'h37B7] = 8'hFF;
DFS[16'h37B8] = 8'hF0;
DFS[16'h37B9] = 8'h6B;
DFS[16'h37BA] = 8'hB1;
DFS[16'h37BB] = 8'hF2;
DFS[16'h37BC] = 8'hC8;
DFS[16'h37BD] = 8'hC9;
DFS[16'h37BE] = 8'h20;
DFS[16'h37BF] = 8'hF0;
DFS[16'h37C0] = 8'hF9;
DFS[16'h37C1] = 8'hB1;
DFS[16'h37C2] = 8'hF2;
DFS[16'h37C3] = 8'h88;
DFS[16'h37C4] = 8'hC9;
DFS[16'h37C5] = 8'h20;
DFS[16'h37C6] = 8'hD0;
DFS[16'h37C7] = 8'h23;
DFS[16'h37C8] = 8'hB1;
DFS[16'h37C9] = 8'hF2;
DFS[16'h37CA] = 8'h38;
DFS[16'h37CB] = 8'hE9;
DFS[16'h37CC] = 8'h30;
DFS[16'h37CD] = 8'h30;
DFS[16'h37CE] = 8'h1C;
DFS[16'h37CF] = 8'hC9;
DFS[16'h37D0] = 8'h0A;
DFS[16'h37D1] = 8'h90;
DFS[16'h37D2] = 8'h14;
DFS[16'h37D3] = 8'hE9;
DFS[16'h37D4] = 8'h07;
DFS[16'h37D5] = 8'hC9;
DFS[16'h37D6] = 8'h0A;
DFS[16'h37D7] = 8'h90;
DFS[16'h37D8] = 8'h12;
DFS[16'h37D9] = 8'hC9;
DFS[16'h37DA] = 8'h10;
DFS[16'h37DB] = 8'h90;
DFS[16'h37DC] = 8'h0A;
DFS[16'h37DD] = 8'hE9;
DFS[16'h37DE] = 8'h20;
DFS[16'h37DF] = 8'hC9;
DFS[16'h37E0] = 8'h0A;
DFS[16'h37E1] = 8'h90;
DFS[16'h37E2] = 8'h08;
DFS[16'h37E3] = 8'hC9;
DFS[16'h37E4] = 8'h10;
DFS[16'h37E5] = 8'hB0;
DFS[16'h37E6] = 8'h04;
DFS[16'h37E7] = 8'hC8;
DFS[16'h37E8] = 8'hC8;
DFS[16'h37E9] = 8'h85;
DFS[16'h37EA] = 8'hA6;
DFS[16'h37EB] = 8'hA5;
DFS[16'h37EC] = 8'hF4;
DFS[16'h37ED] = 8'h85;
DFS[16'h37EE] = 8'hA7;
DFS[16'h37EF] = 8'h98;
DFS[16'h37F0] = 8'h48;
DFS[16'h37F1] = 8'hA0;
DFS[16'h37F2] = 8'h24;
DFS[16'h37F3] = 8'hB9;
DFS[16'h37F4] = 8'hE7;
DFS[16'h37F5] = 8'hB8;
DFS[16'h37F6] = 8'h99;
DFS[16'h37F7] = 8'h52;
DFS[16'h37F8] = 8'h0D;
DFS[16'h37F9] = 8'h88;
DFS[16'h37FA] = 8'h10;
DFS[16'h37FB] = 8'hF7;
DFS[16'h37FC] = 8'hA2;
DFS[16'h37FD] = 8'h0F;
DFS[16'h37FE] = 8'h20;
DFS[16'h37FF] = 8'h52;
DFS[16'h3800] = 8'h0D;
DFS[16'h3801] = 8'h68;
DFS[16'h3802] = 8'hA8;
DFS[16'h3803] = 8'h86;
DFS[16'h3804] = 8'hA6;
DFS[16'h3805] = 8'h8A;
DFS[16'h3806] = 8'h10;
DFS[16'h3807] = 8'h14;
DFS[16'h3808] = 8'h20;
DFS[16'h3809] = 8'h00;
DFS[16'h380A] = 8'hA0;
DFS[16'h380B] = 8'hFF;
DFS[16'h380C] = 8'h4E;
DFS[16'h380D] = 8'h6F;
DFS[16'h380E] = 8'h20;
DFS[16'h380F] = 8'h53;
DFS[16'h3810] = 8'h69;
DFS[16'h3811] = 8'h64;
DFS[16'h3812] = 8'h65;
DFS[16'h3813] = 8'h77;
DFS[16'h3814] = 8'h61;
DFS[16'h3815] = 8'h79;
DFS[16'h3816] = 8'h73;
DFS[16'h3817] = 8'h20;
DFS[16'h3818] = 8'h52;
DFS[16'h3819] = 8'h41;
DFS[16'h381A] = 8'h4D;
DFS[16'h381B] = 8'h00;
DFS[16'h381C] = 8'h20;
DFS[16'h381D] = 8'h62;
DFS[16'h381E] = 8'h82;
DFS[16'h381F] = 8'h18;
DFS[16'h3820] = 8'h20;
DFS[16'h3821] = 8'hC2;
DFS[16'h3822] = 8'hFF;
DFS[16'h3823] = 8'hD0;
DFS[16'h3824] = 8'h03;
DFS[16'h3825] = 8'h4C;
DFS[16'h3826] = 8'hB0;
DFS[16'h3827] = 8'hB2;
DFS[16'h3828] = 8'h20;
DFS[16'h3829] = 8'hFE;
DFS[16'h382A] = 8'h80;
DFS[16'h382B] = 8'h98;
DFS[16'h382C] = 8'h20;
DFS[16'h382D] = 8'h71;
DFS[16'h382E] = 8'h82;
DFS[16'h382F] = 8'hB9;
DFS[16'h3830] = 8'h0E;
DFS[16'h3831] = 8'h0F;
DFS[16'h3832] = 8'h48;
DFS[16'h3833] = 8'h29;
DFS[16'h3834] = 8'h03;
DFS[16'h3835] = 8'h85;
DFS[16'h3836] = 8'hA1;
DFS[16'h3837] = 8'hB9;
DFS[16'h3838] = 8'h0F;
DFS[16'h3839] = 8'h0F;
DFS[16'h383A] = 8'h85;
DFS[16'h383B] = 8'hA0;
DFS[16'h383C] = 8'h68;
DFS[16'h383D] = 8'h4A;
DFS[16'h383E] = 8'h4A;
DFS[16'h383F] = 8'h29;
DFS[16'h3840] = 8'h03;
DFS[16'h3841] = 8'hF0;
DFS[16'h3842] = 8'h04;
DFS[16'h3843] = 8'h49;
DFS[16'h3844] = 8'h03;
DFS[16'h3845] = 8'hD0;
DFS[16'h3846] = 8'h16;
DFS[16'h3847] = 8'hB9;
DFS[16'h3848] = 8'h0C;
DFS[16'h3849] = 8'h0F;
DFS[16'h384A] = 8'hD0;
DFS[16'h384B] = 8'h11;
DFS[16'h384C] = 8'hB9;
DFS[16'h384D] = 8'h0D;
DFS[16'h384E] = 8'h0F;
DFS[16'h384F] = 8'h30;
DFS[16'h3850] = 8'h0C;
DFS[16'h3851] = 8'h85;
DFS[16'h3852] = 8'hA5;
DFS[16'h3853] = 8'hA2;
DFS[16'h3854] = 8'h05;
DFS[16'h3855] = 8'hC9;
DFS[16'h3856] = 8'h40;
DFS[16'h3857] = 8'hF0;
DFS[16'h3858] = 8'h15;
DFS[16'h3859] = 8'h0A;
DFS[16'h385A] = 8'hCA;
DFS[16'h385B] = 8'hD0;
DFS[16'h385C] = 8'hF8;
DFS[16'h385D] = 8'h20;
DFS[16'h385E] = 8'h00;
DFS[16'h385F] = 8'hA0;
DFS[16'h3860] = 8'hFF;
DFS[16'h3861] = 8'h42;
DFS[16'h3862] = 8'h61;
DFS[16'h3863] = 8'h64;
DFS[16'h3864] = 8'h20;
DFS[16'h3865] = 8'h52;
DFS[16'h3866] = 8'h4F;
DFS[16'h3867] = 8'h4D;
DFS[16'h3868] = 8'h20;
DFS[16'h3869] = 8'h73;
DFS[16'h386A] = 8'h69;
DFS[16'h386B] = 8'h7A;
DFS[16'h386C] = 8'h65;
DFS[16'h386D] = 8'h00;
DFS[16'h386E] = 8'h46;
DFS[16'h386F] = 8'hA5;
DFS[16'h3870] = 8'hA6;
DFS[16'h3871] = 8'hCF;
DFS[16'h3872] = 8'h20;
DFS[16'h3873] = 8'h7E;
DFS[16'h3874] = 8'hAA;
DFS[16'h3875] = 8'h18;
DFS[16'h3876] = 8'hA5;
DFS[16'h3877] = 8'hA2;
DFS[16'h3878] = 8'h65;
DFS[16'h3879] = 8'hA0;
DFS[16'h387A] = 8'h85;
DFS[16'h387B] = 8'hA2;
DFS[16'h387C] = 8'hA5;
DFS[16'h387D] = 8'hA3;
DFS[16'h387E] = 8'h65;
DFS[16'h387F] = 8'hA1;
DFS[16'h3880] = 8'h85;
DFS[16'h3881] = 8'hA3;
DFS[16'h3882] = 8'hA9;
DFS[16'h3883] = 8'h00;
DFS[16'h3884] = 8'h65;
DFS[16'h3885] = 8'hA4;
DFS[16'h3886] = 8'h85;
DFS[16'h3887] = 8'hA4;
DFS[16'h3888] = 8'hA0;
DFS[16'h3889] = 8'h1C;
DFS[16'h388A] = 8'hB9;
DFS[16'h388B] = 8'hCB;
DFS[16'h388C] = 8'hB8;
DFS[16'h388D] = 8'h99;
DFS[16'h388E] = 8'h52;
DFS[16'h388F] = 8'h0D;
DFS[16'h3890] = 8'h88;
DFS[16'h3891] = 8'h10;
DFS[16'h3892] = 8'hF7;
DFS[16'h3893] = 8'hA5;
DFS[16'h3894] = 8'hA6;
DFS[16'h3895] = 8'h8D;
DFS[16'h3896] = 8'h53;
DFS[16'h3897] = 8'h0D;
DFS[16'h3898] = 8'hA5;
DFS[16'h3899] = 8'hA7;
DFS[16'h389A] = 8'h8D;
DFS[16'h389B] = 8'h69;
DFS[16'h389C] = 8'h0D;
DFS[16'h389D] = 8'h20;
DFS[16'h389E] = 8'hEC;
DFS[16'h389F] = 8'hA4;
DFS[16'h38A0] = 8'hA9;
DFS[16'h38A1] = 8'hFF;
DFS[16'h38A2] = 8'h8D;
DFS[16'h38A3] = 8'h82;
DFS[16'h38A4] = 8'h10;
DFS[16'h38A5] = 8'h20;
DFS[16'h38A6] = 8'h0F;
DFS[16'h38A7] = 8'hA6;
DFS[16'h38A8] = 8'h20;
DFS[16'h38A9] = 8'h52;
DFS[16'h38AA] = 8'h0D;
DFS[16'h38AB] = 8'h18;
DFS[16'h38AC] = 8'hA5;
DFS[16'h38AD] = 8'hA2;
DFS[16'h38AE] = 8'h69;
DFS[16'h38AF] = 8'h02;
DFS[16'h38B0] = 8'h85;
DFS[16'h38B1] = 8'hA2;
DFS[16'h38B2] = 8'h90;
DFS[16'h38B3] = 8'h06;
DFS[16'h38B4] = 8'hE6;
DFS[16'h38B5] = 8'hA3;
DFS[16'h38B6] = 8'hD0;
DFS[16'h38B7] = 8'h02;
DFS[16'h38B8] = 8'hE6;
DFS[16'h38B9] = 8'hA3;
DFS[16'h38BA] = 8'hEE;
DFS[16'h38BB] = 8'h5E;
DFS[16'h38BC] = 8'h0D;
DFS[16'h38BD] = 8'hEE;
DFS[16'h38BE] = 8'h5E;
DFS[16'h38BF] = 8'h0D;
DFS[16'h38C0] = 8'hEE;
DFS[16'h38C1] = 8'h64;
DFS[16'h38C2] = 8'h0D;
DFS[16'h38C3] = 8'hEE;
DFS[16'h38C4] = 8'h64;
DFS[16'h38C5] = 8'h0D;
DFS[16'h38C6] = 8'hC6;
DFS[16'h38C7] = 8'hA5;
DFS[16'h38C8] = 8'hD0;
DFS[16'h38C9] = 8'hDB;
DFS[16'h38CA] = 8'h60;
DFS[16'h38CB] = 8'hA9;
DFS[16'h38CC] = 8'h00;
DFS[16'h38CD] = 8'h8D;
DFS[16'h38CE] = 8'h30;
DFS[16'h38CF] = 8'hFE;
DFS[16'h38D0] = 8'hA0;
DFS[16'h38D1] = 8'h00;
DFS[16'h38D2] = 8'hB9;
DFS[16'h38D3] = 8'h00;
DFS[16'h38D4] = 8'h0E;
DFS[16'h38D5] = 8'h99;
DFS[16'h38D6] = 8'h00;
DFS[16'h38D7] = 8'h80;
DFS[16'h38D8] = 8'hB9;
DFS[16'h38D9] = 8'h00;
DFS[16'h38DA] = 8'h0F;
DFS[16'h38DB] = 8'h99;
DFS[16'h38DC] = 8'h00;
DFS[16'h38DD] = 8'h81;
DFS[16'h38DE] = 8'h88;
DFS[16'h38DF] = 8'hD0;
DFS[16'h38E0] = 8'hF1;
DFS[16'h38E1] = 8'hA9;
DFS[16'h38E2] = 8'h00;
DFS[16'h38E3] = 8'h8D;
DFS[16'h38E4] = 8'h30;
DFS[16'h38E5] = 8'hFE;
DFS[16'h38E6] = 8'h60;
DFS[16'h38E7] = 8'h8E;
DFS[16'h38E8] = 8'h30;
DFS[16'h38E9] = 8'hFE;
DFS[16'h38EA] = 8'hAD;
DFS[16'h38EB] = 8'hFF;
DFS[16'h38EC] = 8'hBF;
DFS[16'h38ED] = 8'hA8;
DFS[16'h38EE] = 8'h49;
DFS[16'h38EF] = 8'hFF;
DFS[16'h38F0] = 8'h8D;
DFS[16'h38F1] = 8'hFF;
DFS[16'h38F2] = 8'hBF;
DFS[16'h38F3] = 8'h98;
DFS[16'h38F4] = 8'h4D;
DFS[16'h38F5] = 8'hFF;
DFS[16'h38F6] = 8'hBF;
DFS[16'h38F7] = 8'h8C;
DFS[16'h38F8] = 8'hFF;
DFS[16'h38F9] = 8'hBF;
DFS[16'h38FA] = 8'hC9;
DFS[16'h38FB] = 8'hFF;
DFS[16'h38FC] = 8'hD0;
DFS[16'h38FD] = 8'h04;
DFS[16'h38FE] = 8'hC6;
DFS[16'h38FF] = 8'hA6;
DFS[16'h3900] = 8'h30;
DFS[16'h3901] = 8'h03;
DFS[16'h3902] = 8'hCA;
DFS[16'h3903] = 8'h10;
DFS[16'h3904] = 8'hE2;
DFS[16'h3905] = 8'hA5;
DFS[16'h3906] = 8'hA7;
DFS[16'h3907] = 8'h8D;
DFS[16'h3908] = 8'h30;
DFS[16'h3909] = 8'hFE;
DFS[16'h390A] = 8'h60;
DFS[16'h390B] = 8'h48;
DFS[16'h390C] = 8'hA5;
DFS[16'h390D] = 8'hCF;
DFS[16'h390E] = 8'h8D;
DFS[16'h390F] = 8'h20;
DFS[16'h3910] = 8'h0D;
DFS[16'h3911] = 8'h68;
DFS[16'h3912] = 8'h60;
DFS[16'h3913] = 8'hA0;
DFS[16'h3914] = 8'h00;
DFS[16'h3915] = 8'hB1;
DFS[16'h3916] = 8'hB0;
DFS[16'h3917] = 8'h30;
DFS[16'h3918] = 8'h07;
DFS[16'h3919] = 8'h29;
DFS[16'h391A] = 8'h03;
DFS[16'h391B] = 8'h85;
DFS[16'h391C] = 8'hCF;
DFS[16'h391D] = 8'h8D;
DFS[16'h391E] = 8'h20;
DFS[16'h391F] = 8'h0D;
DFS[16'h3920] = 8'hA0;
DFS[16'h3921] = 8'h05;
DFS[16'h3922] = 8'hB1;
DFS[16'h3923] = 8'hB0;
DFS[16'h3924] = 8'h18;
DFS[16'h3925] = 8'h69;
DFS[16'h3926] = 8'h07;
DFS[16'h3927] = 8'h85;
DFS[16'h3928] = 8'hBE;
DFS[16'h3929] = 8'h20;
DFS[16'h392A] = 8'h37;
DFS[16'h392B] = 8'hB9;
DFS[16'h392C] = 8'hA4;
DFS[16'h392D] = 8'hBE;
DFS[16'h392E] = 8'hB0;
DFS[16'h392F] = 8'h02;
DFS[16'h3930] = 8'hA9;
DFS[16'h3931] = 8'h00;
DFS[16'h3932] = 8'h91;
DFS[16'h3933] = 8'hB0;
DFS[16'h3934] = 8'hA9;
DFS[16'h3935] = 8'h00;
DFS[16'h3936] = 8'h60;
DFS[16'h3937] = 8'hC8;
DFS[16'h3938] = 8'hB1;
DFS[16'h3939] = 8'hB0;
DFS[16'h393A] = 8'hAA;
DFS[16'h393B] = 8'h29;
DFS[16'h393C] = 8'h3F;
DFS[16'h393D] = 8'h85;
DFS[16'h393E] = 8'hBF;
DFS[16'h393F] = 8'hC9;
DFS[16'h3940] = 8'h3A;
DFS[16'h3941] = 8'hD0;
DFS[16'h3942] = 8'h2B;
DFS[16'h3943] = 8'hA5;
DFS[16'h3944] = 8'hBE;
DFS[16'h3945] = 8'hC9;
DFS[16'h3946] = 8'h09;
DFS[16'h3947] = 8'hD0;
DFS[16'h3948] = 8'h13;
DFS[16'h3949] = 8'hC8;
DFS[16'h394A] = 8'hB1;
DFS[16'h394B] = 8'hB0;
DFS[16'h394C] = 8'hC9;
DFS[16'h394D] = 8'h23;
DFS[16'h394E] = 8'hD0;
DFS[16'h394F] = 8'h0C;
DFS[16'h3950] = 8'hC8;
DFS[16'h3951] = 8'hB1;
DFS[16'h3952] = 8'hB0;
DFS[16'h3953] = 8'h29;
DFS[16'h3954] = 8'h20;
DFS[16'h3955] = 8'hF0;
DFS[16'h3956] = 8'h02;
DFS[16'h3957] = 8'hA9;
DFS[16'h3958] = 8'h02;
DFS[16'h3959] = 8'h8D;
DFS[16'h395A] = 8'h20;
DFS[16'h395B] = 8'h0D;
DFS[16'h395C] = 8'h18;
DFS[16'h395D] = 8'h60;
DFS[16'h395E] = 8'hA9;
DFS[16'h395F] = 8'h1E;
DFS[16'h3960] = 8'h38;
DFS[16'h3961] = 8'h60;
DFS[16'h3962] = 8'hA9;
DFS[16'h3963] = 8'h10;
DFS[16'h3964] = 8'h38;
DFS[16'h3965] = 8'h60;
DFS[16'h3966] = 8'hA9;
DFS[16'h3967] = 8'h12;
DFS[16'h3968] = 8'h38;
DFS[16'h3969] = 8'h60;
DFS[16'h396A] = 8'hA9;
DFS[16'h396B] = 8'hFF;
DFS[16'h396C] = 8'h38;
DFS[16'h396D] = 8'h60;
DFS[16'h396E] = 8'hA5;
DFS[16'h396F] = 8'hCF;
DFS[16'h3970] = 8'h6A;
DFS[16'h3971] = 8'h8A;
DFS[16'h3972] = 8'h90;
DFS[16'h3973] = 8'h02;
DFS[16'h3974] = 8'h49;
DFS[16'h3975] = 8'hC0;
DFS[16'h3976] = 8'h2A;
DFS[16'h3977] = 8'h90;
DFS[16'h3978] = 8'h0C;
DFS[16'h3979] = 8'h2A;
DFS[16'h397A] = 8'hB0;
DFS[16'h397B] = 8'hE2;
DFS[16'h397C] = 8'hAD;
DFS[16'h397D] = 8'h20;
DFS[16'h397E] = 8'h0D;
DFS[16'h397F] = 8'h29;
DFS[16'h3980] = 8'h02;
DFS[16'h3981] = 8'h09;
DFS[16'h3982] = 8'h01;
DFS[16'h3983] = 8'hD0;
DFS[16'h3984] = 8'h08;
DFS[16'h3985] = 8'h2A;
DFS[16'h3986] = 8'h90;
DFS[16'h3987] = 8'hDA;
DFS[16'h3988] = 8'hAD;
DFS[16'h3989] = 8'h20;
DFS[16'h398A] = 8'h0D;
DFS[16'h398B] = 8'h29;
DFS[16'h398C] = 8'h02;
DFS[16'h398D] = 8'h8D;
DFS[16'h398E] = 8'h20;
DFS[16'h398F] = 8'h0D;
DFS[16'h3990] = 8'hAA;
DFS[16'h3991] = 8'h86;
DFS[16'h3992] = 8'hC0;
DFS[16'h3993] = 8'hBD;
DFS[16'h3994] = 8'h10;
DFS[16'h3995] = 8'h0D;
DFS[16'h3996] = 8'h30;
DFS[16'h3997] = 8'hCA;
DFS[16'h3998] = 8'hA5;
DFS[16'h3999] = 8'hBF;
DFS[16'h399A] = 8'hC9;
DFS[16'h399B] = 8'h13;
DFS[16'h399C] = 8'hF0;
DFS[16'h399D] = 8'h0B;
DFS[16'h399E] = 8'hC9;
DFS[16'h399F] = 8'h0B;
DFS[16'h39A0] = 8'hD0;
DFS[16'h39A1] = 8'hBA;
DFS[16'h39A2] = 8'hBD;
DFS[16'h39A3] = 8'h1C;
DFS[16'h39A4] = 8'h0D;
DFS[16'h39A5] = 8'hC9;
DFS[16'h39A6] = 8'h54;
DFS[16'h39A7] = 8'hD0;
DFS[16'h39A8] = 8'hBD;
DFS[16'h39A9] = 8'hA5;
DFS[16'h39AA] = 8'hBE;
DFS[16'h39AB] = 8'hC9;
DFS[16'h39AC] = 8'h0A;
DFS[16'h39AD] = 8'hD0;
DFS[16'h39AE] = 8'hBB;
DFS[16'h39AF] = 8'h20;
DFS[16'h39B0] = 8'hEC;
DFS[16'h39B1] = 8'hA4;
DFS[16'h39B2] = 8'hA9;
DFS[16'h39B3] = 8'h00;
DFS[16'h39B4] = 8'h85;
DFS[16'h39B5] = 8'hC5;
DFS[16'h39B6] = 8'hC8;
DFS[16'h39B7] = 8'hB1;
DFS[16'h39B8] = 8'hB0;
DFS[16'h39B9] = 8'hC9;
DFS[16'h39BA] = 8'h50;
DFS[16'h39BB] = 8'hB0;
DFS[16'h39BC] = 8'hA1;
DFS[16'h39BD] = 8'h0A;
DFS[16'h39BE] = 8'h85;
DFS[16'h39BF] = 8'hC4;
DFS[16'h39C0] = 8'h0A;
DFS[16'h39C1] = 8'h26;
DFS[16'h39C2] = 8'hC5;
DFS[16'h39C3] = 8'h0A;
DFS[16'h39C4] = 8'h26;
DFS[16'h39C5] = 8'hC5;
DFS[16'h39C6] = 8'h65;
DFS[16'h39C7] = 8'hC4;
DFS[16'h39C8] = 8'h85;
DFS[16'h39C9] = 8'hC4;
DFS[16'h39CA] = 8'h90;
DFS[16'h39CB] = 8'h02;
DFS[16'h39CC] = 8'hE6;
DFS[16'h39CD] = 8'hC5;
DFS[16'h39CE] = 8'hC8;
DFS[16'h39CF] = 8'hB1;
DFS[16'h39D0] = 8'hB0;
DFS[16'h39D1] = 8'hC9;
DFS[16'h39D2] = 8'h0A;
DFS[16'h39D3] = 8'hB0;
DFS[16'h39D4] = 8'h62;
DFS[16'h39D5] = 8'h18;
DFS[16'h39D6] = 8'h65;
DFS[16'h39D7] = 8'hC4;
DFS[16'h39D8] = 8'h85;
DFS[16'h39D9] = 8'hC4;
DFS[16'h39DA] = 8'h90;
DFS[16'h39DB] = 8'h02;
DFS[16'h39DC] = 8'hE6;
DFS[16'h39DD] = 8'hC5;
DFS[16'h39DE] = 8'hC8;
DFS[16'h39DF] = 8'hB1;
DFS[16'h39E0] = 8'hB0;
DFS[16'h39E1] = 8'h29;
DFS[16'h39E2] = 8'h1F;
DFS[16'h39E3] = 8'h85;
DFS[16'h39E4] = 8'hA5;
DFS[16'h39E5] = 8'hF0;
DFS[16'h39E6] = 8'h46;
DFS[16'h39E7] = 8'h18;
DFS[16'h39E8] = 8'h65;
DFS[16'h39E9] = 8'hC4;
DFS[16'h39EA] = 8'hAA;
DFS[16'h39EB] = 8'hA9;
DFS[16'h39EC] = 8'h00;
DFS[16'h39ED] = 8'h65;
DFS[16'h39EE] = 8'hC5;
DFS[16'h39EF] = 8'hC9;
DFS[16'h39F0] = 8'h03;
DFS[16'h39F1] = 8'h90;
DFS[16'h39F2] = 8'h06;
DFS[16'h39F3] = 8'hD0;
DFS[16'h39F4] = 8'h42;
DFS[16'h39F5] = 8'hE0;
DFS[16'h39F6] = 8'h21;
DFS[16'h39F7] = 8'hB0;
DFS[16'h39F8] = 8'h3E;
DFS[16'h39F9] = 8'hA6;
DFS[16'h39FA] = 8'hC0;
DFS[16'h39FB] = 8'hBD;
DFS[16'h39FC] = 8'h10;
DFS[16'h39FD] = 8'h0D;
DFS[16'h39FE] = 8'h6A;
DFS[16'h39FF] = 8'hBD;
DFS[16'h3A00] = 8'h0C;
DFS[16'h3A01] = 8'h0D;
DFS[16'h3A02] = 8'h20;
DFS[16'h3A03] = 8'h87;
DFS[16'h3A04] = 8'hAA;
DFS[16'h3A05] = 8'h18;
DFS[16'h3A06] = 8'hA5;
DFS[16'h3A07] = 8'hA2;
DFS[16'h3A08] = 8'h65;
DFS[16'h3A09] = 8'hC4;
DFS[16'h3A0A] = 8'h85;
DFS[16'h3A0B] = 8'hA2;
DFS[16'h3A0C] = 8'hA5;
DFS[16'h3A0D] = 8'hA3;
DFS[16'h3A0E] = 8'h65;
DFS[16'h3A0F] = 8'hC5;
DFS[16'h3A10] = 8'h85;
DFS[16'h3A11] = 8'hA3;
DFS[16'h3A12] = 8'h90;
DFS[16'h3A13] = 8'h02;
DFS[16'h3A14] = 8'hE6;
DFS[16'h3A15] = 8'hA4;
DFS[16'h3A16] = 8'hA0;
DFS[16'h3A17] = 8'h00;
DFS[16'h3A18] = 8'h84;
DFS[16'h3A19] = 8'hA7;
DFS[16'h3A1A] = 8'hC8;
DFS[16'h3A1B] = 8'hB1;
DFS[16'h3A1C] = 8'hB0;
DFS[16'h3A1D] = 8'h85;
DFS[16'h3A1E] = 8'hA0;
DFS[16'h3A1F] = 8'hC8;
DFS[16'h3A20] = 8'hB1;
DFS[16'h3A21] = 8'hB0;
DFS[16'h3A22] = 8'h85;
DFS[16'h3A23] = 8'hA1;
DFS[16'h3A24] = 8'hA5;
DFS[16'h3A25] = 8'hBF;
DFS[16'h3A26] = 8'hC9;
DFS[16'h3A27] = 8'h13;
DFS[16'h3A28] = 8'hF0;
DFS[16'h3A29] = 8'h05;
DFS[16'h3A2A] = 8'h20;
DFS[16'h3A2B] = 8'hAB;
DFS[16'h3A2C] = 8'hAB;
DFS[16'h3A2D] = 8'h18;
DFS[16'h3A2E] = 8'h60;
DFS[16'h3A2F] = 8'h20;
DFS[16'h3A30] = 8'h42;
DFS[16'h3A31] = 8'hA6;
DFS[16'h3A32] = 8'h20;
DFS[16'h3A33] = 8'hCD;
DFS[16'h3A34] = 8'hA0;
DFS[16'h3A35] = 8'h18;
DFS[16'h3A36] = 8'h60;
DFS[16'h3A37] = 8'hA9;
DFS[16'h3A38] = 8'h1E;
DFS[16'h3A39] = 8'h38;
DFS[16'h3A3A] = 8'h60;
DFS[16'h3A3B] = 8'h54;
DFS[16'h3A3C] = 8'h45;
DFS[16'h3A3D] = 8'h53;
DFS[16'h3A3E] = 8'h53;
DFS[16'h3A3F] = 8'h20;
DFS[16'h3A40] = 8'h54;
DFS[16'h3A41] = 8'h45;
DFS[16'h3A42] = 8'h53;
DFS[16'h3A43] = 8'h53;
DFS[16'h3A44] = 8'h20;
DFS[16'h3A45] = 8'h54;
DFS[16'h3A46] = 8'h45;
DFS[16'h3A47] = 8'h53;
DFS[16'h3A48] = 8'h53;
DFS[16'h3A49] = 8'h20;
DFS[16'h3A4A] = 8'h54;
DFS[16'h3A4B] = 8'h45;
DFS[16'h3A4C] = 8'h53;
DFS[16'h3A4D] = 8'h53;
DFS[16'h3A4E] = 8'h20;
DFS[16'h3A4F] = 8'h54;
DFS[16'h3A50] = 8'h45;
DFS[16'h3A51] = 8'h53;
DFS[16'h3A52] = 8'h53;
DFS[16'h3A53] = 8'h20;
DFS[16'h3A54] = 8'h54;
DFS[16'h3A55] = 8'h45;
DFS[16'h3A56] = 8'h53;
DFS[16'h3A57] = 8'h53;
DFS[16'h3A58] = 8'h20;
DFS[16'h3A59] = 8'h54;
DFS[16'h3A5A] = 8'h45;
DFS[16'h3A5B] = 8'h53;
DFS[16'h3A5C] = 8'h53;
DFS[16'h3A5D] = 8'h20;
DFS[16'h3A5E] = 8'h54;
DFS[16'h3A5F] = 8'h45;
DFS[16'h3A60] = 8'h53;
DFS[16'h3A61] = 8'h53;
DFS[16'h3A62] = 8'h20;
DFS[16'h3A63] = 8'h54;
DFS[16'h3A64] = 8'h45;
DFS[16'h3A65] = 8'h53;
DFS[16'h3A66] = 8'h53;
DFS[16'h3A67] = 8'h20;
DFS[16'h3A68] = 8'h54;
DFS[16'h3A69] = 8'h45;
DFS[16'h3A6A] = 8'h53;
DFS[16'h3A6B] = 8'h53;
DFS[16'h3A6C] = 8'h20;
DFS[16'h3A6D] = 8'h54;
DFS[16'h3A6E] = 8'h45;
DFS[16'h3A6F] = 8'h53;
DFS[16'h3A70] = 8'h53;
DFS[16'h3A71] = 8'h20;
DFS[16'h3A72] = 8'h54;
DFS[16'h3A73] = 8'h45;
DFS[16'h3A74] = 8'h53;
DFS[16'h3A75] = 8'h53;
DFS[16'h3A76] = 8'h20;
DFS[16'h3A77] = 8'h54;
DFS[16'h3A78] = 8'h45;
DFS[16'h3A79] = 8'h53;
DFS[16'h3A7A] = 8'h53;
DFS[16'h3A7B] = 8'h20;
DFS[16'h3A7C] = 8'h54;
DFS[16'h3A7D] = 8'h45;
DFS[16'h3A7E] = 8'h53;
DFS[16'h3A7F] = 8'h53;
DFS[16'h3A80] = 8'h20;
DFS[16'h3A81] = 8'h54;
DFS[16'h3A82] = 8'h45;
DFS[16'h3A83] = 8'h53;
DFS[16'h3A84] = 8'h53;
DFS[16'h3A85] = 8'h20;
DFS[16'h3A86] = 8'h54;
DFS[16'h3A87] = 8'h45;
DFS[16'h3A88] = 8'h53;
DFS[16'h3A89] = 8'h53;
DFS[16'h3A8A] = 8'h20;
DFS[16'h3A8B] = 8'h54;
DFS[16'h3A8C] = 8'h45;
DFS[16'h3A8D] = 8'h53;
DFS[16'h3A8E] = 8'h53;
DFS[16'h3A8F] = 8'h20;
DFS[16'h3A90] = 8'h54;
DFS[16'h3A91] = 8'h45;
DFS[16'h3A92] = 8'h53;
DFS[16'h3A93] = 8'h53;
DFS[16'h3A94] = 8'h20;
DFS[16'h3A95] = 8'h54;
DFS[16'h3A96] = 8'h45;
DFS[16'h3A97] = 8'h53;
DFS[16'h3A98] = 8'h53;
DFS[16'h3A99] = 8'h20;
DFS[16'h3A9A] = 8'h54;
DFS[16'h3A9B] = 8'h45;
DFS[16'h3A9C] = 8'h53;
DFS[16'h3A9D] = 8'h53;
DFS[16'h3A9E] = 8'h20;
DFS[16'h3A9F] = 8'h54;
DFS[16'h3AA0] = 8'h45;
DFS[16'h3AA1] = 8'h53;
DFS[16'h3AA2] = 8'h53;
DFS[16'h3AA3] = 8'h20;
DFS[16'h3AA4] = 8'h54;
DFS[16'h3AA5] = 8'h45;
DFS[16'h3AA6] = 8'h53;
DFS[16'h3AA7] = 8'h53;
DFS[16'h3AA8] = 8'h20;
DFS[16'h3AA9] = 8'h54;
DFS[16'h3AAA] = 8'h45;
DFS[16'h3AAB] = 8'h53;
DFS[16'h3AAC] = 8'h53;
DFS[16'h3AAD] = 8'h20;
DFS[16'h3AAE] = 8'h54;
DFS[16'h3AAF] = 8'h45;
DFS[16'h3AB0] = 8'h53;
DFS[16'h3AB1] = 8'h53;
DFS[16'h3AB2] = 8'h20;
DFS[16'h3AB3] = 8'h54;
DFS[16'h3AB4] = 8'h45;
DFS[16'h3AB5] = 8'h53;
DFS[16'h3AB6] = 8'h53;
DFS[16'h3AB7] = 8'h20;
DFS[16'h3AB8] = 8'h54;
DFS[16'h3AB9] = 8'h45;
DFS[16'h3ABA] = 8'h53;
DFS[16'h3ABB] = 8'h53;
DFS[16'h3ABC] = 8'h20;
DFS[16'h3ABD] = 8'h54;
DFS[16'h3ABE] = 8'h45;
DFS[16'h3ABF] = 8'h53;
DFS[16'h3AC0] = 8'h53;
DFS[16'h3AC1] = 8'h20;
DFS[16'h3AC2] = 8'h54;
DFS[16'h3AC3] = 8'h45;
DFS[16'h3AC4] = 8'h53;
DFS[16'h3AC5] = 8'h53;
DFS[16'h3AC6] = 8'h20;
DFS[16'h3AC7] = 8'h54;
DFS[16'h3AC8] = 8'h45;
DFS[16'h3AC9] = 8'h53;
DFS[16'h3ACA] = 8'h53;
DFS[16'h3ACB] = 8'h20;
DFS[16'h3ACC] = 8'h54;
DFS[16'h3ACD] = 8'h45;
DFS[16'h3ACE] = 8'h53;
DFS[16'h3ACF] = 8'h53;
DFS[16'h3AD0] = 8'h20;
DFS[16'h3AD1] = 8'h54;
DFS[16'h3AD2] = 8'h45;
DFS[16'h3AD3] = 8'h53;
DFS[16'h3AD4] = 8'h53;
DFS[16'h3AD5] = 8'h20;
DFS[16'h3AD6] = 8'h54;
DFS[16'h3AD7] = 8'h45;
DFS[16'h3AD8] = 8'h53;
DFS[16'h3AD9] = 8'h53;
DFS[16'h3ADA] = 8'h20;
DFS[16'h3ADB] = 8'h54;
DFS[16'h3ADC] = 8'h45;
DFS[16'h3ADD] = 8'h53;
DFS[16'h3ADE] = 8'h53;
DFS[16'h3ADF] = 8'h20;
DFS[16'h3AE0] = 8'h54;
DFS[16'h3AE1] = 8'h45;
DFS[16'h3AE2] = 8'h53;
DFS[16'h3AE3] = 8'h53;
DFS[16'h3AE4] = 8'h20;
DFS[16'h3AE5] = 8'h54;
DFS[16'h3AE6] = 8'h45;
DFS[16'h3AE7] = 8'h53;
DFS[16'h3AE8] = 8'h53;
DFS[16'h3AE9] = 8'h20;
DFS[16'h3AEA] = 8'h54;
DFS[16'h3AEB] = 8'h45;
DFS[16'h3AEC] = 8'h53;
DFS[16'h3AED] = 8'h53;
DFS[16'h3AEE] = 8'h20;
DFS[16'h3AEF] = 8'h54;
DFS[16'h3AF0] = 8'h45;
DFS[16'h3AF1] = 8'h53;
DFS[16'h3AF2] = 8'h53;
DFS[16'h3AF3] = 8'h20;
DFS[16'h3AF4] = 8'h54;
DFS[16'h3AF5] = 8'h45;
DFS[16'h3AF6] = 8'h53;
DFS[16'h3AF7] = 8'h53;
DFS[16'h3AF8] = 8'h20;
DFS[16'h3AF9] = 8'h54;
DFS[16'h3AFA] = 8'h45;
DFS[16'h3AFB] = 8'h53;
DFS[16'h3AFC] = 8'h53;
DFS[16'h3AFD] = 8'h20;
DFS[16'h3AFE] = 8'h54;
DFS[16'h3AFF] = 8'h45;
DFS[16'h3B00] = 8'h53;
DFS[16'h3B01] = 8'h53;
DFS[16'h3B02] = 8'h20;
DFS[16'h3B03] = 8'h54;
DFS[16'h3B04] = 8'h45;
DFS[16'h3B05] = 8'h53;
DFS[16'h3B06] = 8'h53;
DFS[16'h3B07] = 8'h20;
DFS[16'h3B08] = 8'h54;
DFS[16'h3B09] = 8'h45;
DFS[16'h3B0A] = 8'h53;
DFS[16'h3B0B] = 8'h53;
DFS[16'h3B0C] = 8'h20;
DFS[16'h3B0D] = 8'h54;
DFS[16'h3B0E] = 8'h45;
DFS[16'h3B0F] = 8'h53;
DFS[16'h3B10] = 8'h53;
DFS[16'h3B11] = 8'h20;
DFS[16'h3B12] = 8'h54;
DFS[16'h3B13] = 8'h45;
DFS[16'h3B14] = 8'h53;
DFS[16'h3B15] = 8'h53;
DFS[16'h3B16] = 8'h20;
DFS[16'h3B17] = 8'h54;
DFS[16'h3B18] = 8'h45;
DFS[16'h3B19] = 8'h53;
DFS[16'h3B1A] = 8'h53;
DFS[16'h3B1B] = 8'h20;
DFS[16'h3B1C] = 8'h54;
DFS[16'h3B1D] = 8'h45;
DFS[16'h3B1E] = 8'h53;
DFS[16'h3B1F] = 8'h53;
DFS[16'h3B20] = 8'h20;
DFS[16'h3B21] = 8'h54;
DFS[16'h3B22] = 8'h45;
DFS[16'h3B23] = 8'h53;
DFS[16'h3B24] = 8'h53;
DFS[16'h3B25] = 8'h20;
DFS[16'h3B26] = 8'h54;
DFS[16'h3B27] = 8'h45;
DFS[16'h3B28] = 8'h53;
DFS[16'h3B29] = 8'h53;
DFS[16'h3B2A] = 8'h20;
DFS[16'h3B2B] = 8'h54;
DFS[16'h3B2C] = 8'h45;
DFS[16'h3B2D] = 8'h53;
DFS[16'h3B2E] = 8'h53;
DFS[16'h3B2F] = 8'h20;
DFS[16'h3B30] = 8'h54;
DFS[16'h3B31] = 8'h45;
DFS[16'h3B32] = 8'h53;
DFS[16'h3B33] = 8'h53;
DFS[16'h3B34] = 8'h20;
DFS[16'h3B35] = 8'h54;
DFS[16'h3B36] = 8'h45;
DFS[16'h3B37] = 8'h53;
DFS[16'h3B38] = 8'h53;
DFS[16'h3B39] = 8'h20;
DFS[16'h3B3A] = 8'h54;
DFS[16'h3B3B] = 8'h45;
DFS[16'h3B3C] = 8'h53;
DFS[16'h3B3D] = 8'h53;
DFS[16'h3B3E] = 8'h20;
DFS[16'h3B3F] = 8'h54;
DFS[16'h3B40] = 8'h45;
DFS[16'h3B41] = 8'h53;
DFS[16'h3B42] = 8'h53;
DFS[16'h3B43] = 8'h20;
DFS[16'h3B44] = 8'h54;
DFS[16'h3B45] = 8'h45;
DFS[16'h3B46] = 8'h53;
DFS[16'h3B47] = 8'h53;
DFS[16'h3B48] = 8'h20;
DFS[16'h3B49] = 8'h54;
DFS[16'h3B4A] = 8'h45;
DFS[16'h3B4B] = 8'h53;
DFS[16'h3B4C] = 8'h53;
DFS[16'h3B4D] = 8'h20;
DFS[16'h3B4E] = 8'h54;
DFS[16'h3B4F] = 8'h45;
DFS[16'h3B50] = 8'h53;
DFS[16'h3B51] = 8'h53;
DFS[16'h3B52] = 8'h20;
DFS[16'h3B53] = 8'h54;
DFS[16'h3B54] = 8'h45;
DFS[16'h3B55] = 8'h53;
DFS[16'h3B56] = 8'h53;
DFS[16'h3B57] = 8'h20;
DFS[16'h3B58] = 8'h54;
DFS[16'h3B59] = 8'h45;
DFS[16'h3B5A] = 8'h53;
DFS[16'h3B5B] = 8'h53;
DFS[16'h3B5C] = 8'h20;
DFS[16'h3B5D] = 8'h54;
DFS[16'h3B5E] = 8'h45;
DFS[16'h3B5F] = 8'h53;
DFS[16'h3B60] = 8'h53;
DFS[16'h3B61] = 8'h20;
DFS[16'h3B62] = 8'h54;
DFS[16'h3B63] = 8'h45;
DFS[16'h3B64] = 8'h53;
DFS[16'h3B65] = 8'h53;
DFS[16'h3B66] = 8'h20;
DFS[16'h3B67] = 8'h54;
DFS[16'h3B68] = 8'h45;
DFS[16'h3B69] = 8'h53;
DFS[16'h3B6A] = 8'h53;
DFS[16'h3B6B] = 8'h20;
DFS[16'h3B6C] = 8'h54;
DFS[16'h3B6D] = 8'h45;
DFS[16'h3B6E] = 8'h53;
DFS[16'h3B6F] = 8'h53;
DFS[16'h3B70] = 8'h20;
DFS[16'h3B71] = 8'h54;
DFS[16'h3B72] = 8'h45;
DFS[16'h3B73] = 8'h53;
DFS[16'h3B74] = 8'h53;
DFS[16'h3B75] = 8'h20;
DFS[16'h3B76] = 8'h54;
DFS[16'h3B77] = 8'h45;
DFS[16'h3B78] = 8'h53;
DFS[16'h3B79] = 8'h53;
DFS[16'h3B7A] = 8'h20;
DFS[16'h3B7B] = 8'h54;
DFS[16'h3B7C] = 8'h45;
DFS[16'h3B7D] = 8'h53;
DFS[16'h3B7E] = 8'h53;
DFS[16'h3B7F] = 8'h20;
DFS[16'h3B80] = 8'h54;
DFS[16'h3B81] = 8'h45;
DFS[16'h3B82] = 8'h53;
DFS[16'h3B83] = 8'h53;
DFS[16'h3B84] = 8'h20;
DFS[16'h3B85] = 8'h54;
DFS[16'h3B86] = 8'h45;
DFS[16'h3B87] = 8'h53;
DFS[16'h3B88] = 8'h53;
DFS[16'h3B89] = 8'h20;
DFS[16'h3B8A] = 8'h54;
DFS[16'h3B8B] = 8'h45;
DFS[16'h3B8C] = 8'h53;
DFS[16'h3B8D] = 8'h53;
DFS[16'h3B8E] = 8'h20;
DFS[16'h3B8F] = 8'h54;
DFS[16'h3B90] = 8'h45;
DFS[16'h3B91] = 8'h53;
DFS[16'h3B92] = 8'h53;
DFS[16'h3B93] = 8'h20;
DFS[16'h3B94] = 8'h54;
DFS[16'h3B95] = 8'h45;
DFS[16'h3B96] = 8'h53;
DFS[16'h3B97] = 8'h53;
DFS[16'h3B98] = 8'h20;
DFS[16'h3B99] = 8'h54;
DFS[16'h3B9A] = 8'h45;
DFS[16'h3B9B] = 8'h53;
DFS[16'h3B9C] = 8'h53;
DFS[16'h3B9D] = 8'h20;
DFS[16'h3B9E] = 8'h54;
DFS[16'h3B9F] = 8'h45;
DFS[16'h3BA0] = 8'h53;
DFS[16'h3BA1] = 8'h53;
DFS[16'h3BA2] = 8'h20;
DFS[16'h3BA3] = 8'h54;
DFS[16'h3BA4] = 8'h45;
DFS[16'h3BA5] = 8'h53;
DFS[16'h3BA6] = 8'h53;
DFS[16'h3BA7] = 8'h20;
DFS[16'h3BA8] = 8'h54;
DFS[16'h3BA9] = 8'h45;
DFS[16'h3BAA] = 8'h53;
DFS[16'h3BAB] = 8'h53;
DFS[16'h3BAC] = 8'h20;
DFS[16'h3BAD] = 8'h54;
DFS[16'h3BAE] = 8'h45;
DFS[16'h3BAF] = 8'h53;
DFS[16'h3BB0] = 8'h53;
DFS[16'h3BB1] = 8'h20;
DFS[16'h3BB2] = 8'h54;
DFS[16'h3BB3] = 8'h45;
DFS[16'h3BB4] = 8'h53;
DFS[16'h3BB5] = 8'h53;
DFS[16'h3BB6] = 8'h20;
DFS[16'h3BB7] = 8'h54;
DFS[16'h3BB8] = 8'h45;
DFS[16'h3BB9] = 8'h53;
DFS[16'h3BBA] = 8'h53;
DFS[16'h3BBB] = 8'h20;
DFS[16'h3BBC] = 8'h54;
DFS[16'h3BBD] = 8'h45;
DFS[16'h3BBE] = 8'h53;
DFS[16'h3BBF] = 8'h53;
DFS[16'h3BC0] = 8'h20;
DFS[16'h3BC1] = 8'h54;
DFS[16'h3BC2] = 8'h45;
DFS[16'h3BC3] = 8'h53;
DFS[16'h3BC4] = 8'h53;
DFS[16'h3BC5] = 8'h20;
DFS[16'h3BC6] = 8'h54;
DFS[16'h3BC7] = 8'h45;
DFS[16'h3BC8] = 8'h53;
DFS[16'h3BC9] = 8'h53;
DFS[16'h3BCA] = 8'h20;
DFS[16'h3BCB] = 8'h54;
DFS[16'h3BCC] = 8'h45;
DFS[16'h3BCD] = 8'h53;
DFS[16'h3BCE] = 8'h53;
DFS[16'h3BCF] = 8'h20;
DFS[16'h3BD0] = 8'h54;
DFS[16'h3BD1] = 8'h45;
DFS[16'h3BD2] = 8'h53;
DFS[16'h3BD3] = 8'h53;
DFS[16'h3BD4] = 8'h20;
DFS[16'h3BD5] = 8'h54;
DFS[16'h3BD6] = 8'h45;
DFS[16'h3BD7] = 8'h53;
DFS[16'h3BD8] = 8'h53;
DFS[16'h3BD9] = 8'h20;
DFS[16'h3BDA] = 8'h54;
DFS[16'h3BDB] = 8'h45;
DFS[16'h3BDC] = 8'h53;
DFS[16'h3BDD] = 8'h53;
DFS[16'h3BDE] = 8'h20;
DFS[16'h3BDF] = 8'h54;
DFS[16'h3BE0] = 8'h45;
DFS[16'h3BE1] = 8'h53;
DFS[16'h3BE2] = 8'h53;
DFS[16'h3BE3] = 8'h20;
DFS[16'h3BE4] = 8'h54;
DFS[16'h3BE5] = 8'h45;
DFS[16'h3BE6] = 8'h53;
DFS[16'h3BE7] = 8'h53;
DFS[16'h3BE8] = 8'h20;
DFS[16'h3BE9] = 8'h54;
DFS[16'h3BEA] = 8'h45;
DFS[16'h3BEB] = 8'h53;
DFS[16'h3BEC] = 8'h53;
DFS[16'h3BED] = 8'h20;
DFS[16'h3BEE] = 8'h54;
DFS[16'h3BEF] = 8'h45;
DFS[16'h3BF0] = 8'h53;
DFS[16'h3BF1] = 8'h53;
DFS[16'h3BF2] = 8'h20;
DFS[16'h3BF3] = 8'h54;
DFS[16'h3BF4] = 8'h45;
DFS[16'h3BF5] = 8'h53;
DFS[16'h3BF6] = 8'h53;
DFS[16'h3BF7] = 8'h20;
DFS[16'h3BF8] = 8'h54;
DFS[16'h3BF9] = 8'h45;
DFS[16'h3BFA] = 8'h53;
DFS[16'h3BFB] = 8'h53;
DFS[16'h3BFC] = 8'h20;
DFS[16'h3BFD] = 8'h54;
DFS[16'h3BFE] = 8'h45;
DFS[16'h3BFF] = 8'h53;
DFS[16'h3C00] = 8'h53;
DFS[16'h3C01] = 8'h20;
DFS[16'h3C02] = 8'h54;
DFS[16'h3C03] = 8'h45;
DFS[16'h3C04] = 8'h53;
DFS[16'h3C05] = 8'h53;
DFS[16'h3C06] = 8'h20;
DFS[16'h3C07] = 8'h54;
DFS[16'h3C08] = 8'h45;
DFS[16'h3C09] = 8'h53;
DFS[16'h3C0A] = 8'h53;
DFS[16'h3C0B] = 8'h20;
DFS[16'h3C0C] = 8'h54;
DFS[16'h3C0D] = 8'h45;
DFS[16'h3C0E] = 8'h53;
DFS[16'h3C0F] = 8'h53;
DFS[16'h3C10] = 8'h20;
DFS[16'h3C11] = 8'h54;
DFS[16'h3C12] = 8'h45;
DFS[16'h3C13] = 8'h53;
DFS[16'h3C14] = 8'h53;
DFS[16'h3C15] = 8'h20;
DFS[16'h3C16] = 8'h54;
DFS[16'h3C17] = 8'h45;
DFS[16'h3C18] = 8'h53;
DFS[16'h3C19] = 8'h53;
DFS[16'h3C1A] = 8'h20;
DFS[16'h3C1B] = 8'h54;
DFS[16'h3C1C] = 8'h45;
DFS[16'h3C1D] = 8'h53;
DFS[16'h3C1E] = 8'h53;
DFS[16'h3C1F] = 8'h20;
DFS[16'h3C20] = 8'h54;
DFS[16'h3C21] = 8'h45;
DFS[16'h3C22] = 8'h53;
DFS[16'h3C23] = 8'h53;
DFS[16'h3C24] = 8'h20;
DFS[16'h3C25] = 8'h54;
DFS[16'h3C26] = 8'h45;
DFS[16'h3C27] = 8'h53;
DFS[16'h3C28] = 8'h53;
DFS[16'h3C29] = 8'h20;
DFS[16'h3C2A] = 8'h54;
DFS[16'h3C2B] = 8'h45;
DFS[16'h3C2C] = 8'h53;
DFS[16'h3C2D] = 8'h53;
DFS[16'h3C2E] = 8'h20;
DFS[16'h3C2F] = 8'h54;
DFS[16'h3C30] = 8'h45;
DFS[16'h3C31] = 8'h53;
DFS[16'h3C32] = 8'h53;
DFS[16'h3C33] = 8'h20;
DFS[16'h3C34] = 8'h54;
DFS[16'h3C35] = 8'h45;
DFS[16'h3C36] = 8'h53;
DFS[16'h3C37] = 8'h53;
DFS[16'h3C38] = 8'h20;
DFS[16'h3C39] = 8'h54;
DFS[16'h3C3A] = 8'h45;
DFS[16'h3C3B] = 8'h53;
DFS[16'h3C3C] = 8'h53;
DFS[16'h3C3D] = 8'h20;
DFS[16'h3C3E] = 8'h54;
DFS[16'h3C3F] = 8'h45;
DFS[16'h3C40] = 8'h53;
DFS[16'h3C41] = 8'h53;
DFS[16'h3C42] = 8'h20;
DFS[16'h3C43] = 8'h54;
DFS[16'h3C44] = 8'h45;
DFS[16'h3C45] = 8'h53;
DFS[16'h3C46] = 8'h53;
DFS[16'h3C47] = 8'h20;
DFS[16'h3C48] = 8'h54;
DFS[16'h3C49] = 8'h45;
DFS[16'h3C4A] = 8'h53;
DFS[16'h3C4B] = 8'h53;
DFS[16'h3C4C] = 8'h20;
DFS[16'h3C4D] = 8'h54;
DFS[16'h3C4E] = 8'h45;
DFS[16'h3C4F] = 8'h53;
DFS[16'h3C50] = 8'h53;
DFS[16'h3C51] = 8'h20;
DFS[16'h3C52] = 8'h54;
DFS[16'h3C53] = 8'h45;
DFS[16'h3C54] = 8'h53;
DFS[16'h3C55] = 8'h53;
DFS[16'h3C56] = 8'h20;
DFS[16'h3C57] = 8'h54;
DFS[16'h3C58] = 8'h45;
DFS[16'h3C59] = 8'h53;
DFS[16'h3C5A] = 8'h53;
DFS[16'h3C5B] = 8'h20;
DFS[16'h3C5C] = 8'h54;
DFS[16'h3C5D] = 8'h45;
DFS[16'h3C5E] = 8'h53;
DFS[16'h3C5F] = 8'h53;
DFS[16'h3C60] = 8'h20;
DFS[16'h3C61] = 8'h54;
DFS[16'h3C62] = 8'h45;
DFS[16'h3C63] = 8'h53;
DFS[16'h3C64] = 8'h53;
DFS[16'h3C65] = 8'h20;
DFS[16'h3C66] = 8'h54;
DFS[16'h3C67] = 8'h45;
DFS[16'h3C68] = 8'h53;
DFS[16'h3C69] = 8'h53;
DFS[16'h3C6A] = 8'h20;
DFS[16'h3C6B] = 8'h54;
DFS[16'h3C6C] = 8'h45;
DFS[16'h3C6D] = 8'h53;
DFS[16'h3C6E] = 8'h53;
DFS[16'h3C6F] = 8'h20;
DFS[16'h3C70] = 8'h54;
DFS[16'h3C71] = 8'h45;
DFS[16'h3C72] = 8'h53;
DFS[16'h3C73] = 8'h53;
DFS[16'h3C74] = 8'h20;
DFS[16'h3C75] = 8'h54;
DFS[16'h3C76] = 8'h45;
DFS[16'h3C77] = 8'h53;
DFS[16'h3C78] = 8'h53;
DFS[16'h3C79] = 8'h20;
DFS[16'h3C7A] = 8'h54;
DFS[16'h3C7B] = 8'h45;
DFS[16'h3C7C] = 8'h53;
DFS[16'h3C7D] = 8'h53;
DFS[16'h3C7E] = 8'h20;
DFS[16'h3C7F] = 8'h54;
DFS[16'h3C80] = 8'h45;
DFS[16'h3C81] = 8'h53;
DFS[16'h3C82] = 8'h53;
DFS[16'h3C83] = 8'h20;
DFS[16'h3C84] = 8'h54;
DFS[16'h3C85] = 8'h45;
DFS[16'h3C86] = 8'h53;
DFS[16'h3C87] = 8'h53;
DFS[16'h3C88] = 8'h20;
DFS[16'h3C89] = 8'h54;
DFS[16'h3C8A] = 8'h45;
DFS[16'h3C8B] = 8'h53;
DFS[16'h3C8C] = 8'h53;
DFS[16'h3C8D] = 8'h20;
DFS[16'h3C8E] = 8'h54;
DFS[16'h3C8F] = 8'h45;
DFS[16'h3C90] = 8'h53;
DFS[16'h3C91] = 8'h53;
DFS[16'h3C92] = 8'h20;
DFS[16'h3C93] = 8'h54;
DFS[16'h3C94] = 8'h45;
DFS[16'h3C95] = 8'h53;
DFS[16'h3C96] = 8'h53;
DFS[16'h3C97] = 8'h20;
DFS[16'h3C98] = 8'h54;
DFS[16'h3C99] = 8'h45;
DFS[16'h3C9A] = 8'h53;
DFS[16'h3C9B] = 8'h53;
DFS[16'h3C9C] = 8'h20;
DFS[16'h3C9D] = 8'h54;
DFS[16'h3C9E] = 8'h45;
DFS[16'h3C9F] = 8'h53;
DFS[16'h3CA0] = 8'h53;
DFS[16'h3CA1] = 8'h20;
DFS[16'h3CA2] = 8'h54;
DFS[16'h3CA3] = 8'h45;
DFS[16'h3CA4] = 8'h53;
DFS[16'h3CA5] = 8'h53;
DFS[16'h3CA6] = 8'h20;
DFS[16'h3CA7] = 8'h54;
DFS[16'h3CA8] = 8'h45;
DFS[16'h3CA9] = 8'h53;
DFS[16'h3CAA] = 8'h53;
DFS[16'h3CAB] = 8'h20;
DFS[16'h3CAC] = 8'h54;
DFS[16'h3CAD] = 8'h45;
DFS[16'h3CAE] = 8'h53;
DFS[16'h3CAF] = 8'h53;
DFS[16'h3CB0] = 8'h20;
DFS[16'h3CB1] = 8'h54;
DFS[16'h3CB2] = 8'h45;
DFS[16'h3CB3] = 8'h53;
DFS[16'h3CB4] = 8'h53;
DFS[16'h3CB5] = 8'h20;
DFS[16'h3CB6] = 8'h54;
DFS[16'h3CB7] = 8'h45;
DFS[16'h3CB8] = 8'h53;
DFS[16'h3CB9] = 8'h53;
DFS[16'h3CBA] = 8'h20;
DFS[16'h3CBB] = 8'h54;
DFS[16'h3CBC] = 8'h45;
DFS[16'h3CBD] = 8'h53;
DFS[16'h3CBE] = 8'h53;
DFS[16'h3CBF] = 8'h20;
DFS[16'h3CC0] = 8'h54;
DFS[16'h3CC1] = 8'h45;
DFS[16'h3CC2] = 8'h53;
DFS[16'h3CC3] = 8'h53;
DFS[16'h3CC4] = 8'h20;
DFS[16'h3CC5] = 8'h54;
DFS[16'h3CC6] = 8'h45;
DFS[16'h3CC7] = 8'h53;
DFS[16'h3CC8] = 8'h53;
DFS[16'h3CC9] = 8'h20;
DFS[16'h3CCA] = 8'h54;
DFS[16'h3CCB] = 8'h45;
DFS[16'h3CCC] = 8'h53;
DFS[16'h3CCD] = 8'h53;
DFS[16'h3CCE] = 8'h20;
DFS[16'h3CCF] = 8'h54;
DFS[16'h3CD0] = 8'h45;
DFS[16'h3CD1] = 8'h53;
DFS[16'h3CD2] = 8'h53;
DFS[16'h3CD3] = 8'h20;
DFS[16'h3CD4] = 8'h54;
DFS[16'h3CD5] = 8'h45;
DFS[16'h3CD6] = 8'h53;
DFS[16'h3CD7] = 8'h53;
DFS[16'h3CD8] = 8'h20;
DFS[16'h3CD9] = 8'h54;
DFS[16'h3CDA] = 8'h45;
DFS[16'h3CDB] = 8'h53;
DFS[16'h3CDC] = 8'h53;
DFS[16'h3CDD] = 8'h20;
DFS[16'h3CDE] = 8'h54;
DFS[16'h3CDF] = 8'h45;
DFS[16'h3CE0] = 8'h53;
DFS[16'h3CE1] = 8'h53;
DFS[16'h3CE2] = 8'h20;
DFS[16'h3CE3] = 8'h54;
DFS[16'h3CE4] = 8'h45;
DFS[16'h3CE5] = 8'h53;
DFS[16'h3CE6] = 8'h53;
DFS[16'h3CE7] = 8'h20;
DFS[16'h3CE8] = 8'h54;
DFS[16'h3CE9] = 8'h45;
DFS[16'h3CEA] = 8'h53;
DFS[16'h3CEB] = 8'h53;
DFS[16'h3CEC] = 8'h20;
DFS[16'h3CED] = 8'h54;
DFS[16'h3CEE] = 8'h45;
DFS[16'h3CEF] = 8'h53;
DFS[16'h3CF0] = 8'h53;
DFS[16'h3CF1] = 8'h20;
DFS[16'h3CF2] = 8'h54;
DFS[16'h3CF3] = 8'h45;
DFS[16'h3CF4] = 8'h53;
DFS[16'h3CF5] = 8'h53;
DFS[16'h3CF6] = 8'h20;
DFS[16'h3CF7] = 8'h54;
DFS[16'h3CF8] = 8'h45;
DFS[16'h3CF9] = 8'h53;
DFS[16'h3CFA] = 8'h53;
DFS[16'h3CFB] = 8'h20;
DFS[16'h3CFC] = 8'h54;
DFS[16'h3CFD] = 8'h45;
DFS[16'h3CFE] = 8'h53;
DFS[16'h3CFF] = 8'h53;
DFS[16'h3D00] = 8'h20;
DFS[16'h3D01] = 8'h54;
DFS[16'h3D02] = 8'h45;
DFS[16'h3D03] = 8'h53;
DFS[16'h3D04] = 8'h53;
DFS[16'h3D05] = 8'h20;
DFS[16'h3D06] = 8'h54;
DFS[16'h3D07] = 8'h45;
DFS[16'h3D08] = 8'h53;
DFS[16'h3D09] = 8'h53;
DFS[16'h3D0A] = 8'h20;
DFS[16'h3D0B] = 8'h54;
DFS[16'h3D0C] = 8'h45;
DFS[16'h3D0D] = 8'h53;
DFS[16'h3D0E] = 8'h53;
DFS[16'h3D0F] = 8'h20;
DFS[16'h3D10] = 8'h54;
DFS[16'h3D11] = 8'h45;
DFS[16'h3D12] = 8'h53;
DFS[16'h3D13] = 8'h53;
DFS[16'h3D14] = 8'h20;
DFS[16'h3D15] = 8'h54;
DFS[16'h3D16] = 8'h45;
DFS[16'h3D17] = 8'h53;
DFS[16'h3D18] = 8'h53;
DFS[16'h3D19] = 8'h20;
DFS[16'h3D1A] = 8'h54;
DFS[16'h3D1B] = 8'h45;
DFS[16'h3D1C] = 8'h53;
DFS[16'h3D1D] = 8'h53;
DFS[16'h3D1E] = 8'h20;
DFS[16'h3D1F] = 8'h54;
DFS[16'h3D20] = 8'h45;
DFS[16'h3D21] = 8'h53;
DFS[16'h3D22] = 8'h53;
DFS[16'h3D23] = 8'h20;
DFS[16'h3D24] = 8'h54;
DFS[16'h3D25] = 8'h45;
DFS[16'h3D26] = 8'h53;
DFS[16'h3D27] = 8'h53;
DFS[16'h3D28] = 8'h20;
DFS[16'h3D29] = 8'h54;
DFS[16'h3D2A] = 8'h45;
DFS[16'h3D2B] = 8'h53;
DFS[16'h3D2C] = 8'h53;
DFS[16'h3D2D] = 8'h20;
DFS[16'h3D2E] = 8'h54;
DFS[16'h3D2F] = 8'h45;
DFS[16'h3D30] = 8'h53;
DFS[16'h3D31] = 8'h53;
DFS[16'h3D32] = 8'h20;
DFS[16'h3D33] = 8'h54;
DFS[16'h3D34] = 8'h45;
DFS[16'h3D35] = 8'h53;
DFS[16'h3D36] = 8'h53;
DFS[16'h3D37] = 8'h20;
DFS[16'h3D38] = 8'h54;
DFS[16'h3D39] = 8'h45;
DFS[16'h3D3A] = 8'h53;
DFS[16'h3D3B] = 8'h53;
DFS[16'h3D3C] = 8'h20;
DFS[16'h3D3D] = 8'h54;
DFS[16'h3D3E] = 8'h45;
DFS[16'h3D3F] = 8'h53;
DFS[16'h3D40] = 8'h53;
DFS[16'h3D41] = 8'h20;
DFS[16'h3D42] = 8'h54;
DFS[16'h3D43] = 8'h45;
DFS[16'h3D44] = 8'h53;
DFS[16'h3D45] = 8'h53;
DFS[16'h3D46] = 8'h20;
DFS[16'h3D47] = 8'h54;
DFS[16'h3D48] = 8'h45;
DFS[16'h3D49] = 8'h53;
DFS[16'h3D4A] = 8'h53;
DFS[16'h3D4B] = 8'h20;
DFS[16'h3D4C] = 8'h54;
DFS[16'h3D4D] = 8'h45;
DFS[16'h3D4E] = 8'h53;
DFS[16'h3D4F] = 8'h53;
DFS[16'h3D50] = 8'h20;
DFS[16'h3D51] = 8'h54;
DFS[16'h3D52] = 8'h45;
DFS[16'h3D53] = 8'h53;
DFS[16'h3D54] = 8'h53;
DFS[16'h3D55] = 8'h20;
DFS[16'h3D56] = 8'h54;
DFS[16'h3D57] = 8'h45;
DFS[16'h3D58] = 8'h53;
DFS[16'h3D59] = 8'h53;
DFS[16'h3D5A] = 8'h20;
DFS[16'h3D5B] = 8'h54;
DFS[16'h3D5C] = 8'h45;
DFS[16'h3D5D] = 8'h53;
DFS[16'h3D5E] = 8'h53;
DFS[16'h3D5F] = 8'h20;
DFS[16'h3D60] = 8'h54;
DFS[16'h3D61] = 8'h45;
DFS[16'h3D62] = 8'h53;
DFS[16'h3D63] = 8'h53;
DFS[16'h3D64] = 8'h20;
DFS[16'h3D65] = 8'h54;
DFS[16'h3D66] = 8'h45;
DFS[16'h3D67] = 8'h53;
DFS[16'h3D68] = 8'h53;
DFS[16'h3D69] = 8'h20;
DFS[16'h3D6A] = 8'h54;
DFS[16'h3D6B] = 8'h45;
DFS[16'h3D6C] = 8'h53;
DFS[16'h3D6D] = 8'h53;
DFS[16'h3D6E] = 8'h20;
DFS[16'h3D6F] = 8'h54;
DFS[16'h3D70] = 8'h45;
DFS[16'h3D71] = 8'h53;
DFS[16'h3D72] = 8'h53;
DFS[16'h3D73] = 8'h20;
DFS[16'h3D74] = 8'h54;
DFS[16'h3D75] = 8'h45;
DFS[16'h3D76] = 8'h53;
DFS[16'h3D77] = 8'h53;
DFS[16'h3D78] = 8'h20;
DFS[16'h3D79] = 8'h54;
DFS[16'h3D7A] = 8'h45;
DFS[16'h3D7B] = 8'h53;
DFS[16'h3D7C] = 8'h53;
DFS[16'h3D7D] = 8'h20;
DFS[16'h3D7E] = 8'h54;
DFS[16'h3D7F] = 8'h45;
DFS[16'h3D80] = 8'h53;
DFS[16'h3D81] = 8'h53;
DFS[16'h3D82] = 8'h20;
DFS[16'h3D83] = 8'h54;
DFS[16'h3D84] = 8'h45;
DFS[16'h3D85] = 8'h53;
DFS[16'h3D86] = 8'h53;
DFS[16'h3D87] = 8'h20;
DFS[16'h3D88] = 8'h54;
DFS[16'h3D89] = 8'h45;
DFS[16'h3D8A] = 8'h53;
DFS[16'h3D8B] = 8'h53;
DFS[16'h3D8C] = 8'h20;
DFS[16'h3D8D] = 8'h54;
DFS[16'h3D8E] = 8'h45;
DFS[16'h3D8F] = 8'h53;
DFS[16'h3D90] = 8'h53;
DFS[16'h3D91] = 8'h20;
DFS[16'h3D92] = 8'h54;
DFS[16'h3D93] = 8'h45;
DFS[16'h3D94] = 8'h53;
DFS[16'h3D95] = 8'h53;
DFS[16'h3D96] = 8'h20;
DFS[16'h3D97] = 8'h54;
DFS[16'h3D98] = 8'h45;
DFS[16'h3D99] = 8'h53;
DFS[16'h3D9A] = 8'h53;
DFS[16'h3D9B] = 8'h20;
DFS[16'h3D9C] = 8'h54;
DFS[16'h3D9D] = 8'h45;
DFS[16'h3D9E] = 8'h53;
DFS[16'h3D9F] = 8'h53;
DFS[16'h3DA0] = 8'h20;
DFS[16'h3DA1] = 8'h54;
DFS[16'h3DA2] = 8'h45;
DFS[16'h3DA3] = 8'h53;
DFS[16'h3DA4] = 8'h53;
DFS[16'h3DA5] = 8'h20;
DFS[16'h3DA6] = 8'h54;
DFS[16'h3DA7] = 8'h45;
DFS[16'h3DA8] = 8'h53;
DFS[16'h3DA9] = 8'h53;
DFS[16'h3DAA] = 8'h20;
DFS[16'h3DAB] = 8'h54;
DFS[16'h3DAC] = 8'h45;
DFS[16'h3DAD] = 8'h53;
DFS[16'h3DAE] = 8'h53;
DFS[16'h3DAF] = 8'h20;
DFS[16'h3DB0] = 8'h54;
DFS[16'h3DB1] = 8'h45;
DFS[16'h3DB2] = 8'h53;
DFS[16'h3DB3] = 8'h53;
DFS[16'h3DB4] = 8'h20;
DFS[16'h3DB5] = 8'h54;
DFS[16'h3DB6] = 8'h45;
DFS[16'h3DB7] = 8'h53;
DFS[16'h3DB8] = 8'h53;
DFS[16'h3DB9] = 8'h20;
DFS[16'h3DBA] = 8'h54;
DFS[16'h3DBB] = 8'h45;
DFS[16'h3DBC] = 8'h53;
DFS[16'h3DBD] = 8'h53;
DFS[16'h3DBE] = 8'h20;
DFS[16'h3DBF] = 8'h54;
DFS[16'h3DC0] = 8'h45;
DFS[16'h3DC1] = 8'h53;
DFS[16'h3DC2] = 8'h53;
DFS[16'h3DC3] = 8'h20;
DFS[16'h3DC4] = 8'h54;
DFS[16'h3DC5] = 8'h45;
DFS[16'h3DC6] = 8'h53;
DFS[16'h3DC7] = 8'h53;
DFS[16'h3DC8] = 8'h20;
DFS[16'h3DC9] = 8'h54;
DFS[16'h3DCA] = 8'h45;
DFS[16'h3DCB] = 8'h53;
DFS[16'h3DCC] = 8'h53;
DFS[16'h3DCD] = 8'h20;
DFS[16'h3DCE] = 8'h54;
DFS[16'h3DCF] = 8'h45;
DFS[16'h3DD0] = 8'h53;
DFS[16'h3DD1] = 8'h53;
DFS[16'h3DD2] = 8'h20;
DFS[16'h3DD3] = 8'h54;
DFS[16'h3DD4] = 8'h45;
DFS[16'h3DD5] = 8'h53;
DFS[16'h3DD6] = 8'h53;
DFS[16'h3DD7] = 8'h20;
DFS[16'h3DD8] = 8'h54;
DFS[16'h3DD9] = 8'h45;
DFS[16'h3DDA] = 8'h53;
DFS[16'h3DDB] = 8'h53;
DFS[16'h3DDC] = 8'h20;
DFS[16'h3DDD] = 8'h54;
DFS[16'h3DDE] = 8'h45;
DFS[16'h3DDF] = 8'h53;
DFS[16'h3DE0] = 8'h53;
DFS[16'h3DE1] = 8'h20;
DFS[16'h3DE2] = 8'h54;
DFS[16'h3DE3] = 8'h45;
DFS[16'h3DE4] = 8'h53;
DFS[16'h3DE5] = 8'h53;
DFS[16'h3DE6] = 8'h20;
DFS[16'h3DE7] = 8'h54;
DFS[16'h3DE8] = 8'h45;
DFS[16'h3DE9] = 8'h53;
DFS[16'h3DEA] = 8'h53;
DFS[16'h3DEB] = 8'h20;
DFS[16'h3DEC] = 8'h54;
DFS[16'h3DED] = 8'h45;
DFS[16'h3DEE] = 8'h53;
DFS[16'h3DEF] = 8'h53;
DFS[16'h3DF0] = 8'h20;
DFS[16'h3DF1] = 8'h54;
DFS[16'h3DF2] = 8'h45;
DFS[16'h3DF3] = 8'h53;
DFS[16'h3DF4] = 8'h53;
DFS[16'h3DF5] = 8'h20;
DFS[16'h3DF6] = 8'h54;
DFS[16'h3DF7] = 8'h45;
DFS[16'h3DF8] = 8'h53;
DFS[16'h3DF9] = 8'h53;
DFS[16'h3DFA] = 8'h20;
DFS[16'h3DFB] = 8'h54;
DFS[16'h3DFC] = 8'h45;
DFS[16'h3DFD] = 8'h53;
DFS[16'h3DFE] = 8'h53;
DFS[16'h3DFF] = 8'h20;
DFS[16'h3E00] = 8'h54;
DFS[16'h3E01] = 8'h45;
DFS[16'h3E02] = 8'h53;
DFS[16'h3E03] = 8'h53;
DFS[16'h3E04] = 8'h20;
DFS[16'h3E05] = 8'h54;
DFS[16'h3E06] = 8'h45;
DFS[16'h3E07] = 8'h53;
DFS[16'h3E08] = 8'h53;
DFS[16'h3E09] = 8'h20;
DFS[16'h3E0A] = 8'h54;
DFS[16'h3E0B] = 8'h45;
DFS[16'h3E0C] = 8'h53;
DFS[16'h3E0D] = 8'h53;
DFS[16'h3E0E] = 8'h20;
DFS[16'h3E0F] = 8'h54;
DFS[16'h3E10] = 8'h45;
DFS[16'h3E11] = 8'h53;
DFS[16'h3E12] = 8'h53;
DFS[16'h3E13] = 8'h20;
DFS[16'h3E14] = 8'h54;
DFS[16'h3E15] = 8'h45;
DFS[16'h3E16] = 8'h53;
DFS[16'h3E17] = 8'h53;
DFS[16'h3E18] = 8'h20;
DFS[16'h3E19] = 8'h54;
DFS[16'h3E1A] = 8'h45;
DFS[16'h3E1B] = 8'h53;
DFS[16'h3E1C] = 8'h53;
DFS[16'h3E1D] = 8'h20;
DFS[16'h3E1E] = 8'h54;
DFS[16'h3E1F] = 8'h45;
DFS[16'h3E20] = 8'h53;
DFS[16'h3E21] = 8'h53;
DFS[16'h3E22] = 8'h20;
DFS[16'h3E23] = 8'h54;
DFS[16'h3E24] = 8'h45;
DFS[16'h3E25] = 8'h53;
DFS[16'h3E26] = 8'h53;
DFS[16'h3E27] = 8'h20;
DFS[16'h3E28] = 8'h54;
DFS[16'h3E29] = 8'h45;
DFS[16'h3E2A] = 8'h53;
DFS[16'h3E2B] = 8'h53;
DFS[16'h3E2C] = 8'h20;
DFS[16'h3E2D] = 8'h54;
DFS[16'h3E2E] = 8'h45;
DFS[16'h3E2F] = 8'h53;
DFS[16'h3E30] = 8'h53;
DFS[16'h3E31] = 8'h20;
DFS[16'h3E32] = 8'h54;
DFS[16'h3E33] = 8'h45;
DFS[16'h3E34] = 8'h53;
DFS[16'h3E35] = 8'h53;
DFS[16'h3E36] = 8'h20;
DFS[16'h3E37] = 8'h54;
DFS[16'h3E38] = 8'h45;
DFS[16'h3E39] = 8'h53;
DFS[16'h3E3A] = 8'h53;
DFS[16'h3E3B] = 8'h20;
DFS[16'h3E3C] = 8'h54;
DFS[16'h3E3D] = 8'h45;
DFS[16'h3E3E] = 8'h53;
DFS[16'h3E3F] = 8'h53;
DFS[16'h3E40] = 8'h20;
DFS[16'h3E41] = 8'h54;
DFS[16'h3E42] = 8'h45;
DFS[16'h3E43] = 8'h53;
DFS[16'h3E44] = 8'h53;
DFS[16'h3E45] = 8'h20;
DFS[16'h3E46] = 8'h54;
DFS[16'h3E47] = 8'h45;
DFS[16'h3E48] = 8'h53;
DFS[16'h3E49] = 8'h53;
DFS[16'h3E4A] = 8'h20;
DFS[16'h3E4B] = 8'h54;
DFS[16'h3E4C] = 8'h45;
DFS[16'h3E4D] = 8'h53;
DFS[16'h3E4E] = 8'h53;
DFS[16'h3E4F] = 8'h20;
DFS[16'h3E50] = 8'h54;
DFS[16'h3E51] = 8'h45;
DFS[16'h3E52] = 8'h53;
DFS[16'h3E53] = 8'h53;
DFS[16'h3E54] = 8'h20;
DFS[16'h3E55] = 8'h54;
DFS[16'h3E56] = 8'h45;
DFS[16'h3E57] = 8'h53;
DFS[16'h3E58] = 8'h53;
DFS[16'h3E59] = 8'h20;
DFS[16'h3E5A] = 8'h54;
DFS[16'h3E5B] = 8'h45;
DFS[16'h3E5C] = 8'h53;
DFS[16'h3E5D] = 8'h53;
DFS[16'h3E5E] = 8'h20;
DFS[16'h3E5F] = 8'h54;
DFS[16'h3E60] = 8'h45;
DFS[16'h3E61] = 8'h53;
DFS[16'h3E62] = 8'h53;
DFS[16'h3E63] = 8'h20;
DFS[16'h3E64] = 8'h54;
DFS[16'h3E65] = 8'h45;
DFS[16'h3E66] = 8'h53;
DFS[16'h3E67] = 8'h53;
DFS[16'h3E68] = 8'h20;
DFS[16'h3E69] = 8'h54;
DFS[16'h3E6A] = 8'h45;
DFS[16'h3E6B] = 8'h53;
DFS[16'h3E6C] = 8'h53;
DFS[16'h3E6D] = 8'h20;
DFS[16'h3E6E] = 8'h54;
DFS[16'h3E6F] = 8'h45;
DFS[16'h3E70] = 8'h53;
DFS[16'h3E71] = 8'h53;
DFS[16'h3E72] = 8'h20;
DFS[16'h3E73] = 8'h54;
DFS[16'h3E74] = 8'h45;
DFS[16'h3E75] = 8'h53;
DFS[16'h3E76] = 8'h53;
DFS[16'h3E77] = 8'h20;
DFS[16'h3E78] = 8'h54;
DFS[16'h3E79] = 8'h45;
DFS[16'h3E7A] = 8'h53;
DFS[16'h3E7B] = 8'h53;
DFS[16'h3E7C] = 8'h20;
DFS[16'h3E7D] = 8'h54;
DFS[16'h3E7E] = 8'h45;
DFS[16'h3E7F] = 8'h53;
DFS[16'h3E80] = 8'h53;
DFS[16'h3E81] = 8'h20;
DFS[16'h3E82] = 8'h54;
DFS[16'h3E83] = 8'h45;
DFS[16'h3E84] = 8'h53;
DFS[16'h3E85] = 8'h53;
DFS[16'h3E86] = 8'h20;
DFS[16'h3E87] = 8'h54;
DFS[16'h3E88] = 8'h45;
DFS[16'h3E89] = 8'h53;
DFS[16'h3E8A] = 8'h53;
DFS[16'h3E8B] = 8'h20;
DFS[16'h3E8C] = 8'h54;
DFS[16'h3E8D] = 8'h45;
DFS[16'h3E8E] = 8'h53;
DFS[16'h3E8F] = 8'h53;
DFS[16'h3E90] = 8'h20;
DFS[16'h3E91] = 8'h54;
DFS[16'h3E92] = 8'h45;
DFS[16'h3E93] = 8'h53;
DFS[16'h3E94] = 8'h53;
DFS[16'h3E95] = 8'h20;
DFS[16'h3E96] = 8'h54;
DFS[16'h3E97] = 8'h45;
DFS[16'h3E98] = 8'h53;
DFS[16'h3E99] = 8'h53;
DFS[16'h3E9A] = 8'h20;
DFS[16'h3E9B] = 8'h54;
DFS[16'h3E9C] = 8'h45;
DFS[16'h3E9D] = 8'h53;
DFS[16'h3E9E] = 8'h53;
DFS[16'h3E9F] = 8'h20;
DFS[16'h3EA0] = 8'h54;
DFS[16'h3EA1] = 8'h45;
DFS[16'h3EA2] = 8'h53;
DFS[16'h3EA3] = 8'h53;
DFS[16'h3EA4] = 8'h20;
DFS[16'h3EA5] = 8'h54;
DFS[16'h3EA6] = 8'h45;
DFS[16'h3EA7] = 8'h53;
DFS[16'h3EA8] = 8'h53;
DFS[16'h3EA9] = 8'h20;
DFS[16'h3EAA] = 8'h54;
DFS[16'h3EAB] = 8'h45;
DFS[16'h3EAC] = 8'h53;
DFS[16'h3EAD] = 8'h53;
DFS[16'h3EAE] = 8'h20;
DFS[16'h3EAF] = 8'h54;
DFS[16'h3EB0] = 8'h45;
DFS[16'h3EB1] = 8'h53;
DFS[16'h3EB2] = 8'h53;
DFS[16'h3EB3] = 8'h20;
DFS[16'h3EB4] = 8'h54;
DFS[16'h3EB5] = 8'h45;
DFS[16'h3EB6] = 8'h53;
DFS[16'h3EB7] = 8'h53;
DFS[16'h3EB8] = 8'h20;
DFS[16'h3EB9] = 8'h54;
DFS[16'h3EBA] = 8'h45;
DFS[16'h3EBB] = 8'h53;
DFS[16'h3EBC] = 8'h53;
DFS[16'h3EBD] = 8'h20;
DFS[16'h3EBE] = 8'h54;
DFS[16'h3EBF] = 8'h45;
DFS[16'h3EC0] = 8'h53;
DFS[16'h3EC1] = 8'h53;
DFS[16'h3EC2] = 8'h20;
DFS[16'h3EC3] = 8'h54;
DFS[16'h3EC4] = 8'h45;
DFS[16'h3EC5] = 8'h53;
DFS[16'h3EC6] = 8'h53;
DFS[16'h3EC7] = 8'h20;
DFS[16'h3EC8] = 8'h54;
DFS[16'h3EC9] = 8'h45;
DFS[16'h3ECA] = 8'h53;
DFS[16'h3ECB] = 8'h53;
DFS[16'h3ECC] = 8'h20;
DFS[16'h3ECD] = 8'h54;
DFS[16'h3ECE] = 8'h45;
DFS[16'h3ECF] = 8'h53;
DFS[16'h3ED0] = 8'h53;
DFS[16'h3ED1] = 8'h20;
DFS[16'h3ED2] = 8'h54;
DFS[16'h3ED3] = 8'h45;
DFS[16'h3ED4] = 8'h53;
DFS[16'h3ED5] = 8'h53;
DFS[16'h3ED6] = 8'h20;
DFS[16'h3ED7] = 8'h54;
DFS[16'h3ED8] = 8'h45;
DFS[16'h3ED9] = 8'h53;
DFS[16'h3EDA] = 8'h53;
DFS[16'h3EDB] = 8'h20;
DFS[16'h3EDC] = 8'h54;
DFS[16'h3EDD] = 8'h45;
DFS[16'h3EDE] = 8'h53;
DFS[16'h3EDF] = 8'h53;
DFS[16'h3EE0] = 8'h20;
DFS[16'h3EE1] = 8'h54;
DFS[16'h3EE2] = 8'h45;
DFS[16'h3EE3] = 8'h53;
DFS[16'h3EE4] = 8'h53;
DFS[16'h3EE5] = 8'h20;
DFS[16'h3EE6] = 8'h54;
DFS[16'h3EE7] = 8'h45;
DFS[16'h3EE8] = 8'h53;
DFS[16'h3EE9] = 8'h53;
DFS[16'h3EEA] = 8'h20;
DFS[16'h3EEB] = 8'h54;
DFS[16'h3EEC] = 8'h45;
DFS[16'h3EED] = 8'h53;
DFS[16'h3EEE] = 8'h53;
DFS[16'h3EEF] = 8'h20;
DFS[16'h3EF0] = 8'h54;
DFS[16'h3EF1] = 8'h45;
DFS[16'h3EF2] = 8'h53;
DFS[16'h3EF3] = 8'h53;
DFS[16'h3EF4] = 8'h20;
DFS[16'h3EF5] = 8'h54;
DFS[16'h3EF6] = 8'h45;
DFS[16'h3EF7] = 8'h53;
DFS[16'h3EF8] = 8'h53;
DFS[16'h3EF9] = 8'h20;
DFS[16'h3EFA] = 8'h54;
DFS[16'h3EFB] = 8'h45;
DFS[16'h3EFC] = 8'h53;
DFS[16'h3EFD] = 8'h53;
DFS[16'h3EFE] = 8'h20;
DFS[16'h3EFF] = 8'h54;
DFS[16'h3F00] = 8'h45;
DFS[16'h3F01] = 8'h53;
DFS[16'h3F02] = 8'h53;
DFS[16'h3F03] = 8'h20;
DFS[16'h3F04] = 8'h54;
DFS[16'h3F05] = 8'h45;
DFS[16'h3F06] = 8'h53;
DFS[16'h3F07] = 8'h53;
DFS[16'h3F08] = 8'h20;
DFS[16'h3F09] = 8'h54;
DFS[16'h3F0A] = 8'h45;
DFS[16'h3F0B] = 8'h53;
DFS[16'h3F0C] = 8'h53;
DFS[16'h3F0D] = 8'h20;
DFS[16'h3F0E] = 8'h54;
DFS[16'h3F0F] = 8'h45;
DFS[16'h3F10] = 8'h53;
DFS[16'h3F11] = 8'h53;
DFS[16'h3F12] = 8'h20;
DFS[16'h3F13] = 8'h54;
DFS[16'h3F14] = 8'h45;
DFS[16'h3F15] = 8'h53;
DFS[16'h3F16] = 8'h53;
DFS[16'h3F17] = 8'h20;
DFS[16'h3F18] = 8'h54;
DFS[16'h3F19] = 8'h45;
DFS[16'h3F1A] = 8'h53;
DFS[16'h3F1B] = 8'h53;
DFS[16'h3F1C] = 8'h20;
DFS[16'h3F1D] = 8'h54;
DFS[16'h3F1E] = 8'h45;
DFS[16'h3F1F] = 8'h53;
DFS[16'h3F20] = 8'h53;
DFS[16'h3F21] = 8'h20;
DFS[16'h3F22] = 8'h54;
DFS[16'h3F23] = 8'h45;
DFS[16'h3F24] = 8'h53;
DFS[16'h3F25] = 8'h53;
DFS[16'h3F26] = 8'h20;
DFS[16'h3F27] = 8'h54;
DFS[16'h3F28] = 8'h45;
DFS[16'h3F29] = 8'h53;
DFS[16'h3F2A] = 8'h53;
DFS[16'h3F2B] = 8'h20;
DFS[16'h3F2C] = 8'h54;
DFS[16'h3F2D] = 8'h45;
DFS[16'h3F2E] = 8'h53;
DFS[16'h3F2F] = 8'h53;
DFS[16'h3F30] = 8'h20;
DFS[16'h3F31] = 8'h54;
DFS[16'h3F32] = 8'h45;
DFS[16'h3F33] = 8'h53;
DFS[16'h3F34] = 8'h53;
DFS[16'h3F35] = 8'h20;
DFS[16'h3F36] = 8'h54;
DFS[16'h3F37] = 8'h45;
DFS[16'h3F38] = 8'h53;
DFS[16'h3F39] = 8'h53;
DFS[16'h3F3A] = 8'h20;
DFS[16'h3F3B] = 8'h54;
DFS[16'h3F3C] = 8'h45;
DFS[16'h3F3D] = 8'h53;
DFS[16'h3F3E] = 8'h53;
DFS[16'h3F3F] = 8'h20;
DFS[16'h3F40] = 8'h54;
DFS[16'h3F41] = 8'h45;
DFS[16'h3F42] = 8'h53;
DFS[16'h3F43] = 8'h53;
DFS[16'h3F44] = 8'h20;
DFS[16'h3F45] = 8'h54;
DFS[16'h3F46] = 8'h45;
DFS[16'h3F47] = 8'h53;
DFS[16'h3F48] = 8'h53;
DFS[16'h3F49] = 8'h20;
DFS[16'h3F4A] = 8'h54;
DFS[16'h3F4B] = 8'h45;
DFS[16'h3F4C] = 8'h53;
DFS[16'h3F4D] = 8'h53;
DFS[16'h3F4E] = 8'h20;
DFS[16'h3F4F] = 8'h54;
DFS[16'h3F50] = 8'h45;
DFS[16'h3F51] = 8'h53;
DFS[16'h3F52] = 8'h53;
DFS[16'h3F53] = 8'h20;
DFS[16'h3F54] = 8'h54;
DFS[16'h3F55] = 8'h45;
DFS[16'h3F56] = 8'h53;
DFS[16'h3F57] = 8'h53;
DFS[16'h3F58] = 8'h20;
DFS[16'h3F59] = 8'h54;
DFS[16'h3F5A] = 8'h45;
DFS[16'h3F5B] = 8'h53;
DFS[16'h3F5C] = 8'h53;
DFS[16'h3F5D] = 8'h20;
DFS[16'h3F5E] = 8'h54;
DFS[16'h3F5F] = 8'h45;
DFS[16'h3F60] = 8'h53;
DFS[16'h3F61] = 8'h53;
DFS[16'h3F62] = 8'h20;
DFS[16'h3F63] = 8'h54;
DFS[16'h3F64] = 8'h45;
DFS[16'h3F65] = 8'h53;
DFS[16'h3F66] = 8'h53;
DFS[16'h3F67] = 8'h20;
DFS[16'h3F68] = 8'h54;
DFS[16'h3F69] = 8'h45;
DFS[16'h3F6A] = 8'h53;
DFS[16'h3F6B] = 8'h53;
DFS[16'h3F6C] = 8'h20;
DFS[16'h3F6D] = 8'h54;
DFS[16'h3F6E] = 8'h45;
DFS[16'h3F6F] = 8'h53;
DFS[16'h3F70] = 8'h53;
DFS[16'h3F71] = 8'h20;
DFS[16'h3F72] = 8'h54;
DFS[16'h3F73] = 8'h45;
DFS[16'h3F74] = 8'h53;
DFS[16'h3F75] = 8'h53;
DFS[16'h3F76] = 8'h20;
DFS[16'h3F77] = 8'h54;
DFS[16'h3F78] = 8'h45;
DFS[16'h3F79] = 8'h53;
DFS[16'h3F7A] = 8'h53;
DFS[16'h3F7B] = 8'h20;
DFS[16'h3F7C] = 8'h54;
DFS[16'h3F7D] = 8'h45;
DFS[16'h3F7E] = 8'h53;
DFS[16'h3F7F] = 8'h53;
DFS[16'h3F80] = 8'h20;
DFS[16'h3F81] = 8'h54;
DFS[16'h3F82] = 8'h45;
DFS[16'h3F83] = 8'h53;
DFS[16'h3F84] = 8'h53;
DFS[16'h3F85] = 8'h20;
DFS[16'h3F86] = 8'h54;
DFS[16'h3F87] = 8'h45;
DFS[16'h3F88] = 8'h53;
DFS[16'h3F89] = 8'h53;
DFS[16'h3F8A] = 8'h20;
DFS[16'h3F8B] = 8'h54;
DFS[16'h3F8C] = 8'h45;
DFS[16'h3F8D] = 8'h53;
DFS[16'h3F8E] = 8'h53;
DFS[16'h3F8F] = 8'h20;
DFS[16'h3F90] = 8'h54;
DFS[16'h3F91] = 8'h45;
DFS[16'h3F92] = 8'h53;
DFS[16'h3F93] = 8'h53;
DFS[16'h3F94] = 8'h20;
DFS[16'h3F95] = 8'h54;
DFS[16'h3F96] = 8'h45;
DFS[16'h3F97] = 8'h53;
DFS[16'h3F98] = 8'h53;
DFS[16'h3F99] = 8'h20;
DFS[16'h3F9A] = 8'h54;
DFS[16'h3F9B] = 8'h45;
DFS[16'h3F9C] = 8'h53;
DFS[16'h3F9D] = 8'h53;
DFS[16'h3F9E] = 8'h20;
DFS[16'h3F9F] = 8'h54;
DFS[16'h3FA0] = 8'h45;
DFS[16'h3FA1] = 8'h53;
DFS[16'h3FA2] = 8'h53;
DFS[16'h3FA3] = 8'h20;
DFS[16'h3FA4] = 8'h54;
DFS[16'h3FA5] = 8'h45;
DFS[16'h3FA6] = 8'h53;
DFS[16'h3FA7] = 8'h53;
DFS[16'h3FA8] = 8'h20;
DFS[16'h3FA9] = 8'h54;
DFS[16'h3FAA] = 8'h45;
DFS[16'h3FAB] = 8'h53;
DFS[16'h3FAC] = 8'h53;
DFS[16'h3FAD] = 8'h20;
DFS[16'h3FAE] = 8'h54;
DFS[16'h3FAF] = 8'h45;
DFS[16'h3FB0] = 8'h53;
DFS[16'h3FB1] = 8'h53;
DFS[16'h3FB2] = 8'h20;
DFS[16'h3FB3] = 8'h54;
DFS[16'h3FB4] = 8'h45;
DFS[16'h3FB5] = 8'h53;
DFS[16'h3FB6] = 8'h53;
DFS[16'h3FB7] = 8'h20;
DFS[16'h3FB8] = 8'h54;
DFS[16'h3FB9] = 8'h45;
DFS[16'h3FBA] = 8'h53;
DFS[16'h3FBB] = 8'h53;
DFS[16'h3FBC] = 8'h20;
DFS[16'h3FBD] = 8'h54;
DFS[16'h3FBE] = 8'h45;
DFS[16'h3FBF] = 8'h53;
DFS[16'h3FC0] = 8'h53;
DFS[16'h3FC1] = 8'h20;
DFS[16'h3FC2] = 8'h54;
DFS[16'h3FC3] = 8'h45;
DFS[16'h3FC4] = 8'h53;
DFS[16'h3FC5] = 8'h53;
DFS[16'h3FC6] = 8'h20;
DFS[16'h3FC7] = 8'h54;
DFS[16'h3FC8] = 8'h45;
DFS[16'h3FC9] = 8'h53;
DFS[16'h3FCA] = 8'h53;
DFS[16'h3FCB] = 8'h20;
DFS[16'h3FCC] = 8'h54;
DFS[16'h3FCD] = 8'h45;
DFS[16'h3FCE] = 8'h53;
DFS[16'h3FCF] = 8'h53;
DFS[16'h3FD0] = 8'h20;
DFS[16'h3FD1] = 8'h54;
DFS[16'h3FD2] = 8'h45;
DFS[16'h3FD3] = 8'h53;
DFS[16'h3FD4] = 8'h53;
DFS[16'h3FD5] = 8'h20;
DFS[16'h3FD6] = 8'h54;
DFS[16'h3FD7] = 8'h45;
DFS[16'h3FD8] = 8'h53;
DFS[16'h3FD9] = 8'h53;
DFS[16'h3FDA] = 8'h20;
DFS[16'h3FDB] = 8'h54;
DFS[16'h3FDC] = 8'h45;
DFS[16'h3FDD] = 8'h53;
DFS[16'h3FDE] = 8'h53;
DFS[16'h3FDF] = 8'h20;
DFS[16'h3FE0] = 8'h54;
DFS[16'h3FE1] = 8'h45;
DFS[16'h3FE2] = 8'h53;
DFS[16'h3FE3] = 8'h53;
DFS[16'h3FE4] = 8'h20;
DFS[16'h3FE5] = 8'h54;
DFS[16'h3FE6] = 8'h45;
DFS[16'h3FE7] = 8'h53;
DFS[16'h3FE8] = 8'h53;
DFS[16'h3FE9] = 8'h20;
DFS[16'h3FEA] = 8'h54;
DFS[16'h3FEB] = 8'h45;
DFS[16'h3FEC] = 8'h53;
DFS[16'h3FED] = 8'h53;
DFS[16'h3FEE] = 8'h20;
DFS[16'h3FEF] = 8'h54;
DFS[16'h3FF0] = 8'h45;
DFS[16'h3FF1] = 8'h53;
DFS[16'h3FF2] = 8'h53;
DFS[16'h3FF3] = 8'h20;
DFS[16'h3FF4] = 8'h54;
DFS[16'h3FF5] = 8'h45;
DFS[16'h3FF6] = 8'h53;
DFS[16'h3FF7] = 8'h53;
DFS[16'h3FF8] = 8'h20;
DFS[16'h3FF9] = 8'h54;
DFS[16'h3FFA] = 8'h45;
DFS[16'h3FFB] = 8'h53;
DFS[16'h3FFC] = 8'h53;
DFS[16'h3FFD] = 8'h20;
DFS[16'h3FFE] = 8'h54;
DFS[16'h3FFF] = 8'h45;
end
