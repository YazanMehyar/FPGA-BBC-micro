`include "TOP.vh"

`define H_COUNT_INIT 799
`define H_PULSE		 784
`define H_BACK		 688
`define H_DISPLAY	 640

`define V_COUNT_INIT 524
`define V_PULSE		 515
`define V_BACK		 513
`define V_DISPLAY	 480
`define V_NEW		 400
