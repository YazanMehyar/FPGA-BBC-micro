`ifndef DEBUG_TOOL
`define DEBUG_TOOL
	`define dl0 6'h00
	`define dl1 6'h01
	`define dl2 6'h02
	`define dl3 6'h03
	`define dl4 6'h04
	`define dl5 6'h05
	`define dl6 6'h06
	`define dl7 6'h07

	`define dl8 6'h08
	`define dl9 6'h09
	`define dlA 6'h0A
	`define dlB 6'h0B
	`define dlC 6'h0C
	`define dlD 6'h0D
	`define dlE 6'h0E
	`define dlF 6'h0F

	`define dlG 6'h10
	`define dlH 6'h11
	`define dlI 6'h12
	`define dlJ 6'h13
	`define dlK 6'h14
	`define dlL 6'h15
	`define dlM 6'h16
	`define dlN 6'h17

	`define dlO 6'h18
	`define dlP 6'h19
	`define dlQ 6'h1A
	`define dlR 6'h1B
	`define dlS 6'h1C
	`define dlT 6'h1D
	`define dlU 6'h1E
	`define dlV 6'h1F

	`define dlW 6'h20
	`define dlX 6'h21
	`define dlY 6'h22
	`define dlZ 6'h23

	`define dlSP 6'h38
	`define SYSVIA 1
	`define USRVIA 0
`endif
