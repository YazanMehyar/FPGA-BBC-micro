`include "TOP.vh"

`define H_DISPLAY 2'b00
`define H_FRONT   2'b01
`define H_PULSE   2'b10
`define H_BACK    2'b11

`define H_COUNTER_INIT 8'd49
`define H_FRONT_COUNT  8'd10
`define H_PULSE_COUNT  8'd9
`define H_BACK_COUNT   8'd3

`define V_DISPLAY 2'b00
`define V_FRONT   2'b01
`define V_PULSE   2'b10
`define V_BACK    2'b11

`define V_COUNTER_INIT 523
`define V_FRONT_COUNT   44
`define V_PULSE_COUNT   33
`define V_BACK_COUNT    31
