`define H_COUNT_INIT 655
`define H_PULSE_INIT 95
`define H_BACKPORCH  47

`define V_COUNT_INIT 490
`define V_PULSE_INIT 1
`define V_BACKPORCH  30

`define PIXELS 640
`define LINES  480
